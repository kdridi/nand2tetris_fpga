LIBRARY ieee;
USE ieee.std_logic_1164.ALL;

ENTITY my_mux8way16_testbench IS
END my_mux8way16_testbench;

ARCHITECTURE behavioral OF my_mux8way16_testbench IS
    COMPONENT my_mux8way16
        PORT (
            a, b, c, d, e, f, g, h : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
            sel : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
            o : OUT STD_LOGIC_VECTOR(15 DOWNTO 0)
        );
    END COMPONENT;

    SIGNAL a, b, c, d, e, f, g, h : STD_LOGIC_VECTOR(15 DOWNTO 0);
    SIGNAL sel : STD_LOGIC_VECTOR(2 DOWNTO 0);
    SIGNAL o_actual : STD_LOGIC_VECTOR(15 DOWNTO 0);
    SIGNAL o_expected : STD_LOGIC_VECTOR(15 DOWNTO 0);

    TYPE test_case IS RECORD
        a, b, c, d, e, f, g, h : STD_LOGIC_VECTOR(15 DOWNTO 0);
        sel : STD_LOGIC_VECTOR(2 DOWNTO 0);
        o : STD_LOGIC_VECTOR(15 DOWNTO 0);
    END RECORD;

    TYPE test_case_array IS ARRAY (NATURAL RANGE <>) OF test_case;
    CONSTANT test_cases : test_case_array := (
        -- a, b, c, d, e, f, g, h, sel, o
        (a => "1011111111111110", b => "1110111001011000", c => "1101110001001101", d => "0100101000000011", e => "1001110001001000", f => "1000011111011011", g => "1011010101101000", h => "1101001010101111", sel => "000", o => "1011111111111110"),
        (a => "0011000000110101", b => "1010111101110001", c => "0001110111011110", d => "0011110000011011", e => "0010100111010011", f => "0100110011101110", g => "1000000001001110", h => "1110011100011101", sel => "001", o => "1010111101110001"),
        (a => "1010110001001000", b => "1000000101001111", c => "1000101110010010", d => "0100100001111110", e => "1111000101001100", f => "1101001100100110", g => "1101100101100001", h => "1100110011000111", sel => "010", o => "1000101110010010"),
        (a => "1101011011011010", b => "0110010110000100", c => "1011011110100000", d => "1101110110011101", e => "1001100100111001", f => "1010100101000011", g => "0111110010000100", h => "0101100100110111", sel => "011", o => "1101110110011101"),
        (a => "1001011110011011", b => "0101100011010001", c => "1010001100111010", d => "0011001111100011", e => "1110000010101100", f => "0101100010100011", g => "0000011010010010", h => "0001000011100001", sel => "100", o => "1110000010101100"),
        (a => "0000100000010100", b => "0010010001110000", c => "0100110011111101", d => "0011000111100111", e => "0111000101011111", f => "1100110101001011", g => "0001100100000100", h => "0001110110100111", sel => "101", o => "1100110101001011"),
        (a => "0100111010011011", b => "1010010010010110", c => "0110011000100101", d => "0011111111100111", e => "0111011110111101", f => "0011111110000110", g => "0000110010101111", h => "0100111010010111", sel => "110", o => "0000110010101111"),
        (a => "1010010100001010", b => "1100010001001111", c => "0010110000110100", d => "0011111001000100", e => "0110110110010011", f => "1010100010111000", g => "1001011101111011", h => "0000010100101110", sel => "111", o => "0000010100101110"),
        (a => "0000000110001001", b => "0011101010110110", c => "0011100100010010", d => "1110001000110110", e => "1001001101011001", f => "0011111110100100", g => "1111001100010111", h => "1001101101101101", sel => "000", o => "0000000110001001"),
        (a => "0110010000010101", b => "0100000000010100", c => "1100110101010100", d => "1101010101110100", e => "0000110101100000", f => "1110011001011000", g => "1111001100011011", h => "0101101111111011", sel => "001", o => "0100000000010100"),
        (a => "1000101011101111", b => "0101100101000000", c => "1001101111100010", d => "0000001010101100", e => "1001100011000110", f => "1010100010010001", g => "0101000101000011", h => "0011110111010000", sel => "010", o => "1001101111100010"),
        (a => "0110110011100001", b => "0111110101110111", c => "0111110000010100", d => "1101101001110100", e => "0010011000110000", f => "0001001110010000", g => "1101111110100010", h => "0010011110111001", sel => "011", o => "1101101001110100"),
        (a => "0100111001000110", b => "0001100010110100", c => "0000100111101111", d => "1110000110011111", e => "0101100001011001", f => "1111110100000111", g => "0111110100001100", h => "1011110001101110", sel => "100", o => "0101100001011001"),
        (a => "0011110100011011", b => "0100101001100000", c => "1001000111100010", d => "0100101001111011", e => "0011000010111000", f => "1000010011111101", g => "1010011001110110", h => "1011101110100111", sel => "101", o => "1000010011111101"),
        (a => "1101111000111101", b => "0100001001011001", c => "1011111001010011", d => "0111011100000011", e => "1110101011101010", f => "0000111110010110", g => "1011010011010011", h => "0101011111001011", sel => "110", o => "1011010011010011"),
        (a => "1000110100001110", b => "0011000011101000", c => "0011001000111111", d => "1011001100111110", e => "0100010001111000", f => "0001000111100010", g => "1101101011110111", h => "1001001010111110", sel => "111", o => "1001001010111110")
    );

    FUNCTION slv_to_string (slv : STD_LOGIC_VECTOR) RETURN STRING IS
        VARIABLE str : STRING (slv'length - 1 DOWNTO 1) := (OTHERS => NUL);
    BEGIN
        FOR n IN slv'length - 1 DOWNTO 1 LOOP
            str(n) := STD_LOGIC'image(slv((n - 1)))(2);
        END LOOP;
        RETURN str;
    END FUNCTION;

BEGIN
    bench : my_mux8way16 PORT MAP(a, b, c, d, e, f, g, h, sel, o_actual);

    PROCESS
    BEGIN

        FOR n IN test_cases'RANGE LOOP
            a <= test_cases(n).a;
            b <= test_cases(n).b;
            c <= test_cases(n).c;
            d <= test_cases(n).d;
            e <= test_cases(n).e;
            f <= test_cases(n).f;
            g <= test_cases(n).g;
            h <= test_cases(n).h;
            sel <= test_cases(n).sel;
            o_expected <= test_cases(n).o;

            WAIT FOR 10 ns;

            ASSERT (o_actual = o_expected)
            REPORT "test failed for " &
                "a = " & slv_to_string(a) &
                ", b = " & slv_to_string(b) &
                ", c = " & slv_to_string(c) &
                ", d = " & slv_to_string(d) &
                ", e = " & slv_to_string(e) &
                ", f = " & slv_to_string(f) &
                ", g = " & slv_to_string(g) &
                ", h = " & slv_to_string(h) &
                ", sel = " & slv_to_string(sel) &
                ". expected o = " & slv_to_string(o_expected) &
                ", got " & slv_to_string(o_actual) SEVERITY error;
        END LOOP;
        WAIT;

    END PROCESS;

END behavioral;