LIBRARY ieee;
USE ieee.std_logic_1164.ALL;

ENTITY my_half_adder_testbench IS
END my_half_adder_testbench;

ARCHITECTURE behavioral OF my_half_adder_testbench IS
    COMPONENT my_half_adder
        PORT (
            a, b : IN STD_LOGIC;
            o : OUT STD_LOGIC;
            c : OUT STD_LOGIC
        );
    END COMPONENT;

    SIGNAL a, b : STD_LOGIC;
    SIGNAL o_actual : STD_LOGIC;
    SIGNAL c_actual : STD_LOGIC;
    SIGNAL o_expected : STD_LOGIC;
    SIGNAL c_expected : STD_LOGIC;

    TYPE test_case IS RECORD
        a, b : STD_LOGIC;
        o : STD_LOGIC;
        c : STD_LOGIC;
    END RECORD;

    TYPE test_case_array IS ARRAY (NATURAL RANGE <>) OF test_case;
    CONSTANT test_cases : test_case_array := (
        -- a, b, o, c
        (a => '0', b => '0', o => '0', c => '0'),
        (a => '0', b => '1', o => '1', c => '0'),
        (a => '1', b => '0', o => '1', c => '0'),
        (a => '1', b => '1', o => '0', c => '1')
    );

    FUNCTION slv_to_string (slv : STD_LOGIC_VECTOR) RETURN STRING IS
        VARIABLE str : STRING (slv'length - 1 DOWNTO 1) := (OTHERS => NUL);
    BEGIN
        FOR n IN slv'length - 1 DOWNTO 1 LOOP
            str(n) := STD_LOGIC'image(slv((n - 1)))(2);
        END LOOP;
        RETURN str;
    END FUNCTION;

BEGIN
    bench : my_half_adder PORT MAP(a, b, o_actual, c_actual);

    PROCESS
    BEGIN

    FOR n IN test_cases'RANGE LOOP
        a <= test_cases(n).a;
        b <= test_cases(n).b;
        o_expected <= test_cases(n).o;
        c_expected <= test_cases(n).c;

        WAIT FOR 10 ns;

        ASSERT (o_actual = o_expected AND c_actual = c_expected)
        REPORT "test failed for " &
            "a = " & STD_LOGIC'image(a) &
            ", b = " & STD_LOGIC'image(b) &
            ". expected o = " & STD_LOGIC'image(o_expected) &
            ", got " & STD_LOGIC'image(o_actual) &
            ". expected c = " & STD_LOGIC'image(c_expected) &
            ", got " & STD_LOGIC'image(c_actual) SEVERITY error;
    END LOOP;
    WAIT;

END PROCESS;

END behavioral;