LIBRARY ieee;
USE ieee.std_logic_1164.ALL;

ENTITY my_alu_testbench IS
END my_alu_testbench;

ARCHITECTURE behavioral OF my_alu_testbench IS
    COMPONENT my_alu
        PORT (
            x, y : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
            zx, nx, zy, ny, f, no : IN STD_LOGIC;
            o : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
            zr, ng : OUT STD_LOGIC
        );
    END COMPONENT;

    SIGNAL x, y : STD_LOGIC_VECTOR(15 DOWNTO 0);
    SIGNAL zx, nx, zy, ny, f, no : STD_LOGIC;
    SIGNAL o_actual : STD_LOGIC_VECTOR(15 DOWNTO 0);
    SIGNAL zr_actual, ng_actual : STD_LOGIC;
    SIGNAL o_expected : STD_LOGIC_VECTOR(15 DOWNTO 0);
    SIGNAL zr_expected, ng_expected : STD_LOGIC;

    TYPE test_case IS RECORD
        x, y : STD_LOGIC_VECTOR(15 DOWNTO 0);
        zx, nx, zy, ny, f, no : STD_LOGIC;
        o : STD_LOGIC_VECTOR(15 DOWNTO 0);
        zr, ng : STD_LOGIC;
    END RECORD;

    TYPE test_case_array IS ARRAY (NATURAL RANGE <>) OF test_case;
    CONSTANT test_cases : test_case_array := (
        -- x, y, zx, nx, zy, ny, f, no, o, zr, ng
        (x => "0000000000000000", y => "1111111111111111", zx => '1', nx => '0', zy => '1', ny => '0', f => '1', no => '0', o => "0000000000000000", zr => '1', ng => '0'),
        (x => "0000000000000000", y => "1111111111111111", zx => '1', nx => '1', zy => '1', ny => '1', f => '1', no => '1', o => "0000000000000001", zr => '0', ng => '0'),
        (x => "0000000000000000", y => "1111111111111111", zx => '1', nx => '1', zy => '1', ny => '0', f => '1', no => '0', o => "1111111111111111", zr => '0', ng => '1'),
        (x => "0000000000000000", y => "1111111111111111", zx => '0', nx => '0', zy => '1', ny => '1', f => '0', no => '0', o => "0000000000000000", zr => '1', ng => '0'),
        (x => "0000000000000000", y => "1111111111111111", zx => '1', nx => '1', zy => '0', ny => '0', f => '0', no => '0', o => "1111111111111111", zr => '0', ng => '1'),
        (x => "0000000000000000", y => "1111111111111111", zx => '0', nx => '0', zy => '1', ny => '1', f => '0', no => '1', o => "1111111111111111", zr => '0', ng => '1'),
        (x => "0000000000000000", y => "1111111111111111", zx => '1', nx => '1', zy => '0', ny => '0', f => '0', no => '1', o => "0000000000000000", zr => '1', ng => '0'),
        (x => "0000000000000000", y => "1111111111111111", zx => '0', nx => '0', zy => '1', ny => '1', f => '1', no => '1', o => "0000000000000000", zr => '1', ng => '0'),
        (x => "0000000000000000", y => "1111111111111111", zx => '1', nx => '1', zy => '0', ny => '0', f => '1', no => '1', o => "0000000000000001", zr => '0', ng => '0'),
        (x => "0000000000000000", y => "1111111111111111", zx => '0', nx => '1', zy => '1', ny => '1', f => '1', no => '1', o => "0000000000000001", zr => '0', ng => '0'),
        (x => "0000000000000000", y => "1111111111111111", zx => '1', nx => '1', zy => '0', ny => '1', f => '1', no => '1', o => "0000000000000000", zr => '1', ng => '0'),
        (x => "0000000000000000", y => "1111111111111111", zx => '0', nx => '0', zy => '1', ny => '1', f => '1', no => '0', o => "1111111111111111", zr => '0', ng => '1'),
        (x => "0000000000000000", y => "1111111111111111", zx => '1', nx => '1', zy => '0', ny => '0', f => '1', no => '0', o => "1111111111111110", zr => '0', ng => '1'),
        (x => "0000000000000000", y => "1111111111111111", zx => '0', nx => '0', zy => '0', ny => '0', f => '1', no => '0', o => "1111111111111111", zr => '0', ng => '1'),
        (x => "0000000000000000", y => "1111111111111111", zx => '0', nx => '1', zy => '0', ny => '0', f => '1', no => '1', o => "0000000000000001", zr => '0', ng => '0'),
        (x => "0000000000000000", y => "1111111111111111", zx => '0', nx => '0', zy => '0', ny => '1', f => '1', no => '1', o => "1111111111111111", zr => '0', ng => '1'),
        (x => "0000000000000000", y => "1111111111111111", zx => '0', nx => '0', zy => '0', ny => '0', f => '0', no => '0', o => "0000000000000000", zr => '1', ng => '0'),
        (x => "0000000000000000", y => "1111111111111111", zx => '0', nx => '1', zy => '0', ny => '1', f => '0', no => '1', o => "1111111111111111", zr => '0', ng => '1'),
        (x => "0000000000010001", y => "0000000000000011", zx => '1', nx => '0', zy => '1', ny => '0', f => '1', no => '0', o => "0000000000000000", zr => '1', ng => '0'),
        (x => "0000000000010001", y => "0000000000000011", zx => '1', nx => '1', zy => '1', ny => '1', f => '1', no => '1', o => "0000000000000001", zr => '0', ng => '0'),
        (x => "0000000000010001", y => "0000000000000011", zx => '1', nx => '1', zy => '1', ny => '0', f => '1', no => '0', o => "1111111111111111", zr => '0', ng => '1'),
        (x => "0000000000010001", y => "0000000000000011", zx => '0', nx => '0', zy => '1', ny => '1', f => '0', no => '0', o => "0000000000010001", zr => '0', ng => '0'),
        (x => "0000000000010001", y => "0000000000000011", zx => '1', nx => '1', zy => '0', ny => '0', f => '0', no => '0', o => "0000000000000011", zr => '0', ng => '0'),
        (x => "0000000000010001", y => "0000000000000011", zx => '0', nx => '0', zy => '1', ny => '1', f => '0', no => '1', o => "1111111111101110", zr => '0', ng => '1'),
        (x => "0000000000010001", y => "0000000000000011", zx => '1', nx => '1', zy => '0', ny => '0', f => '0', no => '1', o => "1111111111111100", zr => '0', ng => '1'),
        (x => "0000000000010001", y => "0000000000000011", zx => '0', nx => '0', zy => '1', ny => '1', f => '1', no => '1', o => "1111111111101111", zr => '0', ng => '1'),
        (x => "0000000000010001", y => "0000000000000011", zx => '1', nx => '1', zy => '0', ny => '0', f => '1', no => '1', o => "1111111111111101", zr => '0', ng => '1'),
        (x => "0000000000010001", y => "0000000000000011", zx => '0', nx => '1', zy => '1', ny => '1', f => '1', no => '1', o => "0000000000010010", zr => '0', ng => '0'),
        (x => "0000000000010001", y => "0000000000000011", zx => '1', nx => '1', zy => '0', ny => '1', f => '1', no => '1', o => "0000000000000100", zr => '0', ng => '0'),
        (x => "0000000000010001", y => "0000000000000011", zx => '0', nx => '0', zy => '1', ny => '1', f => '1', no => '0', o => "0000000000010000", zr => '0', ng => '0'),
        (x => "0000000000010001", y => "0000000000000011", zx => '1', nx => '1', zy => '0', ny => '0', f => '1', no => '0', o => "0000000000000010", zr => '0', ng => '0'),
        (x => "0000000000010001", y => "0000000000000011", zx => '0', nx => '0', zy => '0', ny => '0', f => '1', no => '0', o => "0000000000010100", zr => '0', ng => '0'),
        (x => "0000000000010001", y => "0000000000000011", zx => '0', nx => '1', zy => '0', ny => '0', f => '1', no => '1', o => "0000000000001110", zr => '0', ng => '0'),
        (x => "0000000000010001", y => "0000000000000011", zx => '0', nx => '0', zy => '0', ny => '1', f => '1', no => '1', o => "1111111111110010", zr => '0', ng => '1'),
        (x => "0000000000010001", y => "0000000000000011", zx => '0', nx => '0', zy => '0', ny => '0', f => '0', no => '0', o => "0000000000000001", zr => '0', ng => '0'),
        (x => "0000000000010001", y => "0000000000000011", zx => '0', nx => '1', zy => '0', ny => '1', f => '0', no => '1', o => "0000000000010011", zr => '0', ng => '0'),
        -- general test cases
        (x => "1000001010111110", y => "1101000001010101", zx => '1', nx => '1', zy => '0', ny => '1', f => '1', no => '1', o => "1101000001010110", zr => '0', ng => '1'),
        (x => "0111111100011001", y => "1111001011111001", zx => '0', nx => '0', zy => '1', ny => '1', f => '1', no => '1', o => "1000000011100111", zr => '0', ng => '1'),
        (x => "1010010011011100", y => "0011011000100111", zx => '1', nx => '1', zy => '1', ny => '1', f => '0', no => '1', o => "0000000000000000", zr => '1', ng => '0'),
        (x => "1111001000010010", y => "1010111110100011", zx => '1', nx => '0', zy => '0', ny => '1', f => '1', no => '1', o => "1010111110100011", zr => '0', ng => '1'),
        (x => "0101011000001101", y => "0100110110111000", zx => '1', nx => '1', zy => '0', ny => '0', f => '1', no => '0', o => "0100110110110111", zr => '0', ng => '0'),
        (x => "0101001000110110", y => "0010111001010111", zx => '1', nx => '1', zy => '1', ny => '1', f => '1', no => '1', o => "0000000000000001", zr => '0', ng => '0'),
        (x => "0001001110011111", y => "1101101111100111", zx => '1', nx => '1', zy => '1', ny => '1', f => '0', no => '1', o => "0000000000000000", zr => '1', ng => '0'),
        (x => "1000111101000101", y => "0111101010011011", zx => '1', nx => '0', zy => '0', ny => '1', f => '0', no => '0', o => "0000000000000000", zr => '1', ng => '0'),
        (x => "1001011110010000", y => "0111110011001101", zx => '0', nx => '1', zy => '1', ny => '0', f => '1', no => '1', o => "1001011110010000", zr => '0', ng => '1'),
        (x => "1011001010010110", y => "0100101000110000", zx => '1', nx => '1', zy => '1', ny => '0', f => '1', no => '0', o => "1111111111111111", zr => '0', ng => '1'),
        (x => "1000110001101000", y => "0011000011111101", zx => '0', nx => '1', zy => '0', ny => '0', f => '0', no => '0', o => "0011000010010101", zr => '0', ng => '0'),
        (x => "1101111011101001", y => "1001011100111100", zx => '1', nx => '1', zy => '1', ny => '1', f => '0', no => '1', o => "0000000000000000", zr => '1', ng => '0'),
        (x => "0101010111110110", y => "0101000011011101", zx => '1', nx => '1', zy => '1', ny => '1', f => '1', no => '1', o => "0000000000000001", zr => '0', ng => '0'),
        (x => "1101010111100010", y => "1001010110000011", zx => '1', nx => '1', zy => '0', ny => '1', f => '0', no => '1', o => "1001010110000011", zr => '0', ng => '1'),
        (x => "1110100001001011", y => "1001011010111100", zx => '1', nx => '1', zy => '1', ny => '1', f => '1', no => '0', o => "1111111111111110", zr => '0', ng => '1'),
        (x => "1100100111100100", y => "1111101010100011", zx => '1', nx => '1', zy => '1', ny => '0', f => '1', no => '1', o => "0000000000000000", zr => '1', ng => '0'),
        (x => "0011111110100111", y => "0000000000010111", zx => '0', nx => '1', zy => '1', ny => '1', f => '0', no => '1', o => "0011111110100111", zr => '0', ng => '0'),
        (x => "0101000110000110", y => "1110001101000100", zx => '1', nx => '1', zy => '0', ny => '0', f => '1', no => '1', o => "0001110010111100", zr => '0', ng => '0'),
        (x => "0010111011000010", y => "1000111111101100", zx => '0', nx => '1', zy => '0', ny => '0', f => '1', no => '1', o => "1001111011010110", zr => '0', ng => '1'),
        (x => "0000111100111100", y => "1011110011101111", zx => '1', nx => '0', zy => '1', ny => '1', f => '0', no => '0', o => "0000000000000000", zr => '1', ng => '0'),
        (x => "0101101100100011", y => "0110100010010000", zx => '1', nx => '0', zy => '1', ny => '0', f => '0', no => '0', o => "0000000000000000", zr => '1', ng => '0'),
        (x => "0111111111011110", y => "1010011111001100", zx => '0', nx => '1', zy => '1', ny => '0', f => '0', no => '0', o => "0000000000000000", zr => '1', ng => '0'),
        (x => "0000011110001010", y => "0001100100010110", zx => '0', nx => '0', zy => '1', ny => '0', f => '0', no => '1', o => "1111111111111111", zr => '0', ng => '1'),
        (x => "0101100100010001", y => "1000111000000110", zx => '1', nx => '1', zy => '0', ny => '1', f => '1', no => '1', o => "1000111000000111", zr => '0', ng => '1'),
        (x => "1001010101010000", y => "1111000001010000", zx => '1', nx => '0', zy => '0', ny => '0', f => '1', no => '1', o => "0000111110101111", zr => '0', ng => '0'),
        (x => "0001101110000100", y => "0011110110100001", zx => '0', nx => '1', zy => '1', ny => '0', f => '1', no => '1', o => "0001101110000100", zr => '0', ng => '0'),
        (x => "1101110110011100", y => "0110001001001100", zx => '0', nx => '0', zy => '0', ny => '1', f => '1', no => '0', o => "0111101101001111", zr => '0', ng => '0'),
        (x => "0110101110000011", y => "0110100000101000", zx => '1', nx => '1', zy => '1', ny => '1', f => '1', no => '1', o => "0000000000000001", zr => '0', ng => '0'),
        (x => "0011110011000111", y => "1100001111101011", zx => '1', nx => '0', zy => '0', ny => '0', f => '0', no => '0', o => "0000000000000000", zr => '1', ng => '0'),
        (x => "0101000110111001", y => "1111110110110010", zx => '1', nx => '1', zy => '1', ny => '0', f => '0', no => '1', o => "1111111111111111", zr => '0', ng => '1'),
        (x => "1101101010110100", y => "0100101010101010", zx => '0', nx => '0', zy => '1', ny => '0', f => '0', no => '1', o => "1111111111111111", zr => '0', ng => '1'),
        (x => "0101101101111100", y => "1000110011101100", zx => '1', nx => '0', zy => '0', ny => '1', f => '1', no => '1', o => "1000110011101100", zr => '0', ng => '1'),
        (x => "0100010011110110", y => "1111111010111001", zx => '1', nx => '1', zy => '1', ny => '0', f => '0', no => '0', o => "0000000000000000", zr => '1', ng => '0'),
        (x => "1011010000000111", y => "0111111000111111", zx => '0', nx => '0', zy => '0', ny => '0', f => '1', no => '1', o => "1100110110111001", zr => '0', ng => '1'),
        (x => "0111100111110000", y => "1100000100110011", zx => '0', nx => '1', zy => '0', ny => '1', f => '0', no => '1', o => "1111100111110011", zr => '0', ng => '1'),
        (x => "0110100000001010", y => "0001111000000011", zx => '0', nx => '0', zy => '1', ny => '1', f => '1', no => '1', o => "1001011111110110", zr => '0', ng => '1'),
        (x => "0001100110111111", y => "0011011101110001", zx => '0', nx => '1', zy => '0', ny => '1', f => '0', no => '1', o => "0011111111111111", zr => '0', ng => '0'),
        (x => "1010111010011111", y => "1111110010011110", zx => '0', nx => '1', zy => '0', ny => '1', f => '0', no => '0', o => "0000000101100000", zr => '0', ng => '0'),
        (x => "1110111101010110", y => "0010000100011110", zx => '0', nx => '0', zy => '0', ny => '1', f => '1', no => '0', o => "1100111000110111", zr => '0', ng => '1'),
        (x => "1001101110110001", y => "1011010001001010", zx => '0', nx => '0', zy => '1', ny => '1', f => '0', no => '0', o => "1001101110110001", zr => '0', ng => '1'),
        (x => "0011010010111100", y => "0111111101100010", zx => '0', nx => '0', zy => '1', ny => '0', f => '1', no => '0', o => "0011010010111100", zr => '0', ng => '0'),
        (x => "1010001101011010", y => "1101110001011110", zx => '1', nx => '1', zy => '1', ny => '0', f => '1', no => '1', o => "0000000000000000", zr => '1', ng => '0'),
        (x => "1001101101100110", y => "1011110011111111", zx => '0', nx => '1', zy => '1', ny => '0', f => '1', no => '1', o => "1001101101100110", zr => '0', ng => '1'),
        (x => "0000010111100000", y => "1010000110011110", zx => '0', nx => '0', zy => '0', ny => '1', f => '1', no => '0', o => "0110010001000001", zr => '0', ng => '0'),
        (x => "1010111101000101", y => "1101001111100011", zx => '1', nx => '0', zy => '0', ny => '0', f => '0', no => '1', o => "1111111111111111", zr => '0', ng => '1'),
        (x => "1001011011010110", y => "1100000100010001", zx => '1', nx => '0', zy => '0', ny => '1', f => '0', no => '1', o => "1111111111111111", zr => '0', ng => '1'),
        (x => "0001111101001011", y => "0011100011100010", zx => '0', nx => '0', zy => '1', ny => '0', f => '1', no => '0', o => "0001111101001011", zr => '0', ng => '0'),
        (x => "0000101111101011", y => "0100000101111000", zx => '0', nx => '1', zy => '1', ny => '0', f => '0', no => '1', o => "1111111111111111", zr => '0', ng => '1'),
        (x => "1111011110101111", y => "0111010010011111", zx => '1', nx => '1', zy => '1', ny => '0', f => '1', no => '0', o => "1111111111111111", zr => '0', ng => '1'),
        (x => "1111111000100011", y => "0111110110000000", zx => '1', nx => '0', zy => '0', ny => '1', f => '1', no => '0', o => "1000001001111111", zr => '0', ng => '1'),
        (x => "0011101101010100", y => "0111111010011111", zx => '0', nx => '1', zy => '0', ny => '1', f => '0', no => '1', o => "0111111111011111", zr => '0', ng => '0'),
        (x => "1100101011100010", y => "1011101110110000", zx => '0', nx => '0', zy => '1', ny => '1', f => '0', no => '1', o => "0011010100011101", zr => '0', ng => '0'),
        (x => "1001001011000010", y => "1101110010000110", zx => '1', nx => '1', zy => '0', ny => '1', f => '0', no => '1', o => "1101110010000110", zr => '0', ng => '1'),
        (x => "0101011101000011", y => "1110111100001000", zx => '1', nx => '0', zy => '0', ny => '0', f => '0', no => '0', o => "0000000000000000", zr => '1', ng => '0'),
        (x => "1110000000010100", y => "1000111100111001", zx => '0', nx => '0', zy => '0', ny => '0', f => '1', no => '0', o => "0110111101001101", zr => '0', ng => '0'),
        (x => "0000010001110000", y => "0101110110000011", zx => '0', nx => '1', zy => '0', ny => '0', f => '0', no => '0', o => "0101100110000011", zr => '0', ng => '0'),
        (x => "0101100100101000", y => "0000010010010011", zx => '1', nx => '1', zy => '0', ny => '1', f => '0', no => '1', o => "0000010010010011", zr => '0', ng => '0'),
        (x => "0100011100001110", y => "1101101110110100", zx => '0', nx => '1', zy => '0', ny => '1', f => '0', no => '0', o => "0010000001000001", zr => '0', ng => '0'),
        (x => "0011001000001000", y => "0101011111110000", zx => '1', nx => '1', zy => '1', ny => '0', f => '0', no => '0', o => "0000000000000000", zr => '1', ng => '0'),
        (x => "0000000110011000", y => "0100110111110101", zx => '1', nx => '1', zy => '0', ny => '0', f => '0', no => '1', o => "1011001000001010", zr => '0', ng => '1'),
        (x => "0100100010111000", y => "0101101111100110", zx => '1', nx => '0', zy => '0', ny => '1', f => '1', no => '1', o => "0101101111100110", zr => '0', ng => '0'),
        (x => "1111110010101111", y => "1100100101001110", zx => '1', nx => '0', zy => '1', ny => '1', f => '1', no => '1', o => "0000000000000000", zr => '1', ng => '0'),
        (x => "1111000011001000", y => "0011110101010001", zx => '1', nx => '1', zy => '1', ny => '1', f => '0', no => '0', o => "1111111111111111", zr => '0', ng => '1'),
        (x => "0110010011111010", y => "1011111110100110", zx => '1', nx => '1', zy => '0', ny => '1', f => '0', no => '0', o => "0100000001011001", zr => '0', ng => '0'),
        (x => "0100011111001001", y => "1110100111001111", zx => '0', nx => '1', zy => '0', ny => '1', f => '0', no => '0', o => "0001000000110000", zr => '0', ng => '0'),
        (x => "1001100110000111", y => "0010101000110001", zx => '1', nx => '0', zy => '1', ny => '0', f => '0', no => '0', o => "0000000000000000", zr => '1', ng => '0'),
        (x => "1101010110111000", y => "1000110010011110", zx => '0', nx => '0', zy => '0', ny => '0', f => '0', no => '0', o => "1000010010011000", zr => '0', ng => '1'),
        (x => "0011101110001010", y => "1111101001011010", zx => '0', nx => '1', zy => '0', ny => '0', f => '1', no => '0', o => "1011111011001111", zr => '0', ng => '1'),
        (x => "0111010101001101", y => "1111111101101101", zx => '0', nx => '1', zy => '1', ny => '1', f => '1', no => '0', o => "1000101010110001", zr => '0', ng => '1'),
        (x => "0100101010011010", y => "1100100011100101", zx => '1', nx => '1', zy => '1', ny => '1', f => '0', no => '0', o => "1111111111111111", zr => '0', ng => '1'),
        (x => "1001111100111110", y => "0000011010111111", zx => '0', nx => '1', zy => '1', ny => '1', f => '1', no => '1', o => "1001111100111111", zr => '0', ng => '1'),
        (x => "1000001010011011", y => "1000001110101100", zx => '1', nx => '1', zy => '0', ny => '0', f => '0', no => '0', o => "1000001110101100", zr => '0', ng => '1'),
        (x => "1000100011001101", y => "1100000010011000", zx => '1', nx => '1', zy => '1', ny => '0', f => '0', no => '0', o => "0000000000000000", zr => '1', ng => '0'),
        (x => "0101010100001000", y => "0011000001110101", zx => '0', nx => '0', zy => '0', ny => '0', f => '1', no => '0', o => "1000010101111101", zr => '0', ng => '1'),
        (x => "0000000101110100", y => "1101101101111110", zx => '0', nx => '1', zy => '0', ny => '1', f => '0', no => '1', o => "1101101101111110", zr => '0', ng => '1'),
        (x => "1111010001011101", y => "0011111111001010", zx => '0', nx => '0', zy => '0', ny => '1', f => '1', no => '1', o => "0100101101101101", zr => '0', ng => '0'),
        (x => "1010011010101000", y => "1000110010001111", zx => '1', nx => '1', zy => '0', ny => '0', f => '1', no => '1', o => "0111001101110001", zr => '0', ng => '0'),
        (x => "1001110010000000", y => "1110110010000101", zx => '1', nx => '0', zy => '1', ny => '0', f => '1', no => '0', o => "0000000000000000", zr => '1', ng => '0'),
        (x => "1110110011100111", y => "1110011100011011", zx => '1', nx => '0', zy => '1', ny => '0', f => '0', no => '1', o => "1111111111111111", zr => '0', ng => '1'),
        (x => "1110111011010101", y => "1000011000110101", zx => '1', nx => '0', zy => '1', ny => '1', f => '1', no => '1', o => "0000000000000000", zr => '1', ng => '0'),
        (x => "0110010000111111", y => "1011010001011111", zx => '1', nx => '1', zy => '0', ny => '1', f => '1', no => '1', o => "1011010001100000", zr => '0', ng => '1'),
        (x => "0011101001100011", y => "0000111010111011", zx => '1', nx => '0', zy => '1', ny => '0', f => '0', no => '0', o => "0000000000000000", zr => '1', ng => '0'),
        (x => "0100010110000010", y => "0111011100010001", zx => '0', nx => '0', zy => '0', ny => '1', f => '0', no => '0', o => "0000000010000010", zr => '0', ng => '0'),
        (x => "0001101011101010", y => "0011100100101010", zx => '1', nx => '1', zy => '0', ny => '1', f => '1', no => '1', o => "0011100100101011", zr => '0', ng => '0'),
        (x => "1000101101000011", y => "0011010010110110", zx => '0', nx => '1', zy => '0', ny => '0', f => '0', no => '1', o => "1100101101001011", zr => '0', ng => '1'),
        (x => "1110101101110011", y => "0000010100011001", zx => '1', nx => '1', zy => '1', ny => '1', f => '1', no => '0', o => "1111111111111110", zr => '0', ng => '1'),
        (x => "0101111111110001", y => "0111011001011000", zx => '0', nx => '0', zy => '0', ny => '0', f => '0', no => '1', o => "1010100110101111", zr => '0', ng => '1'),
        (x => "0110100011110101", y => "0110011111101110", zx => '1', nx => '1', zy => '1', ny => '1', f => '0', no => '0', o => "1111111111111111", zr => '0', ng => '1'),
        (x => "0111101111111100", y => "1110000011110111", zx => '0', nx => '0', zy => '0', ny => '0', f => '0', no => '0', o => "0110000011110100", zr => '0', ng => '0'),
        (x => "1110001101110110", y => "1001101000011101", zx => '1', nx => '0', zy => '1', ny => '1', f => '0', no => '0', o => "0000000000000000", zr => '1', ng => '0'),
        (x => "0100001110111000", y => "0011011001001011", zx => '1', nx => '1', zy => '0', ny => '1', f => '1', no => '1', o => "0011011001001100", zr => '0', ng => '0'),
        (x => "0110101111101001", y => "0010000111100111", zx => '0', nx => '1', zy => '1', ny => '1', f => '1', no => '0', o => "1001010000010101", zr => '0', ng => '1'),
        (x => "0001100010111110", y => "1110101010010101", zx => '1', nx => '1', zy => '0', ny => '1', f => '1', no => '0', o => "0001010101101001", zr => '0', ng => '0'),
        (x => "0011100101100000", y => "0011010001001011", zx => '1', nx => '1', zy => '0', ny => '0', f => '0', no => '1', o => "1100101110110100", zr => '0', ng => '1'),
        (x => "0001100110100100", y => "0000100001001001", zx => '1', nx => '0', zy => '1', ny => '0', f => '0', no => '1', o => "1111111111111111", zr => '0', ng => '1'),
        (x => "0010101011010000", y => "1001011110100011", zx => '1', nx => '0', zy => '1', ny => '1', f => '1', no => '0', o => "1111111111111111", zr => '0', ng => '1'),
        (x => "1000001001001111", y => "0101110011100100", zx => '1', nx => '0', zy => '1', ny => '0', f => '1', no => '0', o => "0000000000000000", zr => '1', ng => '0'),
        (x => "0111001001110001", y => "1110101100001001", zx => '0', nx => '0', zy => '0', ny => '1', f => '1', no => '0', o => "1000011101100111", zr => '0', ng => '1'),
        (x => "1001100101111010", y => "0100110110101010", zx => '0', nx => '0', zy => '0', ny => '0', f => '0', no => '0', o => "0000100100101010", zr => '0', ng => '0'),
        (x => "0100111000101010", y => "0100000011010011", zx => '1', nx => '0', zy => '0', ny => '0', f => '1', no => '0', o => "0100000011010011", zr => '0', ng => '0'),
        (x => "1110101101101111", y => "1100010001010100", zx => '0', nx => '1', zy => '1', ny => '1', f => '0', no => '0', o => "0001010010010000", zr => '0', ng => '0'),
        (x => "1000100011010011", y => "0000111100000001", zx => '1', nx => '1', zy => '1', ny => '0', f => '1', no => '1', o => "0000000000000000", zr => '1', ng => '0'),
        (x => "1111000000110010", y => "1010011011111011", zx => '1', nx => '1', zy => '1', ny => '0', f => '0', no => '0', o => "0000000000000000", zr => '1', ng => '0'),
        (x => "0011111000101001", y => "1101110110001011", zx => '1', nx => '0', zy => '0', ny => '0', f => '0', no => '0', o => "0000000000000000", zr => '1', ng => '0'),
        (x => "1001001101010010", y => "0001011110110010", zx => '0', nx => '1', zy => '1', ny => '1', f => '1', no => '1', o => "1001001101010011", zr => '0', ng => '1'),
        (x => "0110101100111001", y => "1111001111000001", zx => '0', nx => '1', zy => '1', ny => '1', f => '0', no => '1', o => "0110101100111001", zr => '0', ng => '0'),
        (x => "0111101110111010", y => "0010010010000011", zx => '1', nx => '1', zy => '1', ny => '0', f => '0', no => '0', o => "0000000000000000", zr => '1', ng => '0'),
        (x => "0111001011110110", y => "0100111000101010", zx => '0', nx => '0', zy => '1', ny => '0', f => '0', no => '0', o => "0000000000000000", zr => '1', ng => '0'),
        (x => "1111111111111110", y => "0111010110101100", zx => '1', nx => '1', zy => '1', ny => '0', f => '0', no => '0', o => "0000000000000000", zr => '1', ng => '0'),
        (x => "0100010011000011", y => "1000100101001101", zx => '0', nx => '0', zy => '0', ny => '1', f => '1', no => '0', o => "1011101101110101", zr => '0', ng => '1'),
        (x => "1011001000100101", y => "0010111011001011", zx => '0', nx => '0', zy => '0', ny => '1', f => '0', no => '1', o => "0110111111011011", zr => '0', ng => '0'),
        (x => "1000011000010111", y => "1010101010110111", zx => '1', nx => '1', zy => '1', ny => '1', f => '0', no => '1', o => "0000000000000000", zr => '1', ng => '0'),
        (x => "1100001001110101", y => "1001101000000100", zx => '0', nx => '1', zy => '1', ny => '0', f => '0', no => '0', o => "0000000000000000", zr => '1', ng => '0'),
        (x => "1100010110010000", y => "0001101000000000", zx => '0', nx => '1', zy => '0', ny => '1', f => '0', no => '0', o => "0010000001101111", zr => '0', ng => '0'),
        (x => "1001101100101011", y => "1011000001100110", zx => '0', nx => '0', zy => '1', ny => '0', f => '0', no => '0', o => "0000000000000000", zr => '1', ng => '0'),
        (x => "0000110001111011", y => "1010110011000110", zx => '1', nx => '0', zy => '0', ny => '0', f => '0', no => '1', o => "1111111111111111", zr => '0', ng => '1'),
        (x => "1111111101101100", y => "0111101011111000", zx => '0', nx => '1', zy => '0', ny => '0', f => '0', no => '1', o => "1111111101101111", zr => '0', ng => '1'),
        (x => "0011101111010110", y => "0010010100010001", zx => '0', nx => '1', zy => '0', ny => '1', f => '1', no => '1', o => "0110000011101000", zr => '0', ng => '0'),
        (x => "0100111000110010", y => "0110101100000101", zx => '0', nx => '0', zy => '1', ny => '0', f => '0', no => '1', o => "1111111111111111", zr => '0', ng => '1'),
        (x => "1100111101010001", y => "1011011010011100", zx => '0', nx => '1', zy => '1', ny => '0', f => '1', no => '1', o => "1100111101010001", zr => '0', ng => '1'),
        (x => "0010011000111000", y => "1101010101000110", zx => '1', nx => '0', zy => '0', ny => '1', f => '0', no => '0', o => "0000000000000000", zr => '1', ng => '0'),
        (x => "0100010100101110", y => "1111101010101010", zx => '1', nx => '0', zy => '1', ny => '1', f => '0', no => '0', o => "0000000000000000", zr => '1', ng => '0'),
        (x => "1011111010110001", y => "1000111100110111", zx => '1', nx => '1', zy => '1', ny => '1', f => '1', no => '1', o => "0000000000000001", zr => '0', ng => '0'),
        (x => "0111100010111100", y => "1101110110000001", zx => '0', nx => '1', zy => '1', ny => '0', f => '1', no => '0', o => "1000011101000011", zr => '0', ng => '1'),
        (x => "1010010000100010", y => "1011011000010010", zx => '1', nx => '1', zy => '1', ny => '0', f => '0', no => '1', o => "1111111111111111", zr => '0', ng => '1'),
        (x => "1110000101011001", y => "1110010010011100", zx => '0', nx => '1', zy => '1', ny => '1', f => '1', no => '0', o => "0001111010100101", zr => '0', ng => '0'),
        (x => "1000010001101100", y => "0111110110100110", zx => '1', nx => '1', zy => '0', ny => '0', f => '1', no => '1', o => "1000001001011010", zr => '0', ng => '1'),
        (x => "1100010010110101", y => "0000000100110111", zx => '0', nx => '0', zy => '0', ny => '1', f => '1', no => '0', o => "1100001101111101", zr => '0', ng => '1'),
        (x => "1011001110000100", y => "1000100011011111", zx => '1', nx => '1', zy => '0', ny => '0', f => '1', no => '0', o => "1000100011011110", zr => '0', ng => '1'),
        (x => "1100001000111111", y => "1001011100001011", zx => '1', nx => '1', zy => '0', ny => '1', f => '1', no => '1', o => "1001011100001100", zr => '0', ng => '1'),
        (x => "1010100011010110", y => "0111001111110101", zx => '1', nx => '0', zy => '0', ny => '0', f => '1', no => '0', o => "0111001111110101", zr => '0', ng => '0'),
        (x => "1111111101010101", y => "1110111001100000", zx => '0', nx => '1', zy => '1', ny => '0', f => '0', no => '0', o => "0000000000000000", zr => '1', ng => '0'),
        (x => "1111001010100110", y => "0101001100010000", zx => '0', nx => '1', zy => '0', ny => '0', f => '0', no => '0', o => "0000000100010000", zr => '0', ng => '0'),
        (x => "0110010100100101", y => "0111110111010110", zx => '1', nx => '1', zy => '1', ny => '0', f => '0', no => '1', o => "1111111111111111", zr => '0', ng => '1'),
        (x => "0101001011110001", y => "0100100011101111", zx => '0', nx => '1', zy => '1', ny => '1', f => '1', no => '0', o => "1010110100001101", zr => '0', ng => '1'),
        (x => "1100100111111000", y => "0011101101001111", zx => '1', nx => '1', zy => '0', ny => '1', f => '1', no => '1', o => "0011101101010000", zr => '0', ng => '0'),
        (x => "1010110001110111", y => "0111111000101010", zx => '1', nx => '0', zy => '0', ny => '1', f => '1', no => '0', o => "1000000111010101", zr => '0', ng => '1'),
        (x => "0010101011100110", y => "1011110110011000", zx => '1', nx => '1', zy => '0', ny => '1', f => '1', no => '0', o => "0100001001100110", zr => '0', ng => '0'),
        (x => "1110110111010010", y => "0110000001000010", zx => '0', nx => '0', zy => '0', ny => '1', f => '0', no => '1', o => "0111001001101111", zr => '0', ng => '0'),
        (x => "1010011011101000", y => "1001000100001100", zx => '0', nx => '0', zy => '1', ny => '0', f => '1', no => '1', o => "0101100100010111", zr => '0', ng => '0'),
        (x => "1000111011100111", y => "1101110110101110", zx => '1', nx => '1', zy => '1', ny => '1', f => '1', no => '0', o => "1111111111111110", zr => '0', ng => '1'),
        (x => "0000000111001101", y => "0010111101100011", zx => '1', nx => '1', zy => '0', ny => '1', f => '1', no => '0', o => "1101000010011011", zr => '0', ng => '1'),
        (x => "0000111110011101", y => "0010101110000101", zx => '0', nx => '0', zy => '1', ny => '1', f => '0', no => '0', o => "0000111110011101", zr => '0', ng => '0'),
        (x => "0000001101000110", y => "0000110011100100", zx => '0', nx => '0', zy => '1', ny => '1', f => '1', no => '1', o => "1111110010111010", zr => '0', ng => '1'),
        (x => "0100101101110000", y => "1111100010111100", zx => '0', nx => '0', zy => '0', ny => '0', f => '1', no => '0', o => "0100010000101100", zr => '0', ng => '0'),
        (x => "0100001110101100", y => "0001010101100111", zx => '1', nx => '1', zy => '1', ny => '0', f => '1', no => '0', o => "1111111111111111", zr => '0', ng => '1'),
        (x => "1001011010001010", y => "1101000100000001", zx => '0', nx => '0', zy => '0', ny => '0', f => '1', no => '0', o => "0110011110001011", zr => '0', ng => '0'),
        (x => "0111111000000001", y => "1111010110110101", zx => '0', nx => '0', zy => '1', ny => '0', f => '0', no => '1', o => "1111111111111111", zr => '0', ng => '1'),
        (x => "1011000110011100", y => "1100111111011111", zx => '1', nx => '0', zy => '0', ny => '1', f => '1', no => '1', o => "1100111111011111", zr => '0', ng => '1'),
        (x => "0010011001010011", y => "0000101001101001", zx => '0', nx => '0', zy => '1', ny => '1', f => '0', no => '1', o => "1101100110101100", zr => '0', ng => '1'),
        (x => "1110101011010001", y => "1101111101001010", zx => '1', nx => '1', zy => '1', ny => '1', f => '0', no => '1', o => "0000000000000000", zr => '1', ng => '0'),
        (x => "1001101100000101", y => "1010100011001000", zx => '1', nx => '0', zy => '1', ny => '1', f => '0', no => '0', o => "0000000000000000", zr => '1', ng => '0'),
        (x => "1000001000010101", y => "0011001001111100", zx => '0', nx => '0', zy => '0', ny => '0', f => '0', no => '1', o => "1111110111101011", zr => '0', ng => '1'),
        (x => "0011100110000101", y => "1100110111010110", zx => '1', nx => '1', zy => '1', ny => '0', f => '0', no => '0', o => "0000000000000000", zr => '1', ng => '0'),
        (x => "1111001110010000", y => "1111010010001010", zx => '1', nx => '0', zy => '0', ny => '1', f => '1', no => '1', o => "1111010010001010", zr => '0', ng => '1'),
        (x => "0001110111010111", y => "0111110001101100", zx => '0', nx => '0', zy => '1', ny => '0', f => '1', no => '0', o => "0001110111010111", zr => '0', ng => '0'),
        (x => "0001001100111100", y => "1001010010010111", zx => '1', nx => '0', zy => '0', ny => '0', f => '0', no => '1', o => "1111111111111111", zr => '0', ng => '1'),
        (x => "0111001011011011", y => "0001010100110010", zx => '1', nx => '0', zy => '0', ny => '0', f => '0', no => '1', o => "1111111111111111", zr => '0', ng => '1'),
        (x => "0101101110100001", y => "0010110101111010", zx => '0', nx => '1', zy => '0', ny => '0', f => '0', no => '0', o => "0010010001011010", zr => '0', ng => '0'),
        (x => "1110111111001100", y => "0101110110110101", zx => '1', nx => '1', zy => '0', ny => '0', f => '1', no => '1', o => "1010001001001011", zr => '0', ng => '1'),
        (x => "0110011100111101", y => "1110011000011011", zx => '1', nx => '0', zy => '0', ny => '1', f => '1', no => '1', o => "1110011000011011", zr => '0', ng => '1'),
        (x => "0111110111101000", y => "1101010001010101", zx => '1', nx => '0', zy => '0', ny => '0', f => '0', no => '0', o => "0000000000000000", zr => '1', ng => '0'),
        (x => "1011001011101111", y => "0010010101101000", zx => '0', nx => '0', zy => '0', ny => '1', f => '0', no => '1', o => "0110110101111000", zr => '0', ng => '0'),
        (x => "0001010010010111", y => "0101010110111010", zx => '0', nx => '1', zy => '0', ny => '0', f => '0', no => '0', o => "0100000100101000", zr => '0', ng => '0'),
        (x => "0101110001000100", y => "0100110100010100", zx => '0', nx => '1', zy => '1', ny => '0', f => '0', no => '0', o => "0000000000000000", zr => '1', ng => '0'),
        (x => "1011011100001101", y => "0011110111011111", zx => '1', nx => '0', zy => '0', ny => '0', f => '0', no => '0', o => "0000000000000000", zr => '1', ng => '0'),
        (x => "1100010011100100", y => "0001011000001110", zx => '0', nx => '0', zy => '1', ny => '1', f => '0', no => '0', o => "1100010011100100", zr => '0', ng => '1'),
        (x => "0011011101010000", y => "1000110101000011", zx => '0', nx => '0', zy => '0', ny => '0', f => '0', no => '0', o => "0000010101000000", zr => '0', ng => '0'),
        (x => "0010011001100111", y => "1010100111011100", zx => '1', nx => '0', zy => '0', ny => '1', f => '0', no => '0', o => "0000000000000000", zr => '1', ng => '0'),
        (x => "0110101001010111", y => "1110101011111010", zx => '1', nx => '0', zy => '1', ny => '0', f => '1', no => '0', o => "0000000000000000", zr => '1', ng => '0'),
        (x => "1101010110101101", y => "0110111110101011", zx => '0', nx => '0', zy => '1', ny => '1', f => '0', no => '1', o => "0010101001010010", zr => '0', ng => '0'),
        (x => "0010000010001011", y => "1011100010111001", zx => '0', nx => '0', zy => '1', ny => '0', f => '0', no => '1', o => "1111111111111111", zr => '0', ng => '1'),
        (x => "1000000101101011", y => "1100101010111101", zx => '1', nx => '0', zy => '1', ny => '1', f => '1', no => '1', o => "0000000000000000", zr => '1', ng => '0'),
        (x => "1000111110000110", y => "1000011110111001", zx => '0', nx => '1', zy => '1', ny => '1', f => '1', no => '0', o => "0111000001111000", zr => '0', ng => '0'),
        (x => "1010001011010100", y => "0001011001011111", zx => '0', nx => '1', zy => '1', ny => '0', f => '0', no => '1', o => "1111111111111111", zr => '0', ng => '1'),
        (x => "1111110010000010", y => "0110010011100111", zx => '1', nx => '0', zy => '1', ny => '1', f => '0', no => '1', o => "1111111111111111", zr => '0', ng => '1'),
        (x => "0011110010001110", y => "1101101110101001", zx => '1', nx => '0', zy => '0', ny => '1', f => '1', no => '1', o => "1101101110101001", zr => '0', ng => '1'),
        (x => "1010010100111010", y => "0010010010001010", zx => '1', nx => '1', zy => '0', ny => '1', f => '0', no => '1', o => "0010010010001010", zr => '0', ng => '0'),
        (x => "1010100101110000", y => "1100100100111100", zx => '0', nx => '1', zy => '0', ny => '0', f => '1', no => '1', o => "1110000000110100", zr => '0', ng => '1'),
        (x => "1101000000101001", y => "0000101101110100", zx => '0', nx => '0', zy => '0', ny => '1', f => '0', no => '1', o => "0010111111110110", zr => '0', ng => '0'),
        (x => "1011101011000000", y => "1001011001100100", zx => '0', nx => '0', zy => '0', ny => '1', f => '0', no => '1', o => "1101011101111111", zr => '0', ng => '1'),
        (x => "1010011101110010", y => "0111010001101011", zx => '0', nx => '1', zy => '1', ny => '1', f => '1', no => '1', o => "1010011101110011", zr => '0', ng => '1'),
        (x => "0001100010000110", y => "1110100001000111", zx => '1', nx => '0', zy => '1', ny => '1', f => '0', no => '1', o => "1111111111111111", zr => '0', ng => '1'),
        (x => "0010110011000011", y => "1100011100100110", zx => '1', nx => '1', zy => '1', ny => '0', f => '1', no => '0', o => "1111111111111111", zr => '0', ng => '1'),
        (x => "1001000100111000", y => "0101000101110011", zx => '1', nx => '1', zy => '0', ny => '1', f => '0', no => '1', o => "0101000101110011", zr => '0', ng => '0'),
        (x => "0101101100010001", y => "1110001111101101", zx => '0', nx => '1', zy => '0', ny => '0', f => '0', no => '0', o => "1010000011101100", zr => '0', ng => '1'),
        (x => "0101110011100101", y => "0001011101111110", zx => '1', nx => '1', zy => '1', ny => '1', f => '0', no => '1', o => "0000000000000000", zr => '1', ng => '0'),
        (x => "0110011101111111", y => "0000010001110001", zx => '0', nx => '1', zy => '1', ny => '1', f => '1', no => '0', o => "1001100001111111", zr => '0', ng => '1'),
        (x => "1100010011100110", y => "0000101010101110", zx => '1', nx => '1', zy => '0', ny => '1', f => '0', no => '0', o => "1111010101010001", zr => '0', ng => '1'),
        (x => "0101011111000011", y => "1001000000000011", zx => '1', nx => '1', zy => '0', ny => '1', f => '1', no => '0', o => "0110111111111011", zr => '0', ng => '0'),
        (x => "1101100111101010", y => "0100100000000000", zx => '0', nx => '1', zy => '1', ny => '0', f => '1', no => '0', o => "0010011000010101", zr => '0', ng => '0'),
        (x => "1110101010000101", y => "1000011111011111", zx => '0', nx => '0', zy => '0', ny => '0', f => '1', no => '1', o => "1000110110011011", zr => '0', ng => '1'),
        (x => "1101011011111110", y => "0100111111100001", zx => '1', nx => '0', zy => '1', ny => '0', f => '1', no => '1', o => "1111111111111111", zr => '0', ng => '1'),
        (x => "1111111010001110", y => "1100001110101010", zx => '1', nx => '1', zy => '1', ny => '1', f => '1', no => '1', o => "0000000000000001", zr => '0', ng => '0'),
        (x => "1100010100101111", y => "0111011010101011", zx => '0', nx => '1', zy => '1', ny => '1', f => '1', no => '0', o => "0011101011001111", zr => '0', ng => '0'),
        (x => "0111001011011101", y => "0101101011110110", zx => '0', nx => '0', zy => '1', ny => '0', f => '0', no => '1', o => "1111111111111111", zr => '0', ng => '1'),
        (x => "1111101100111001", y => "1000011111100100", zx => '0', nx => '0', zy => '0', ny => '1', f => '0', no => '0', o => "0111100000011001", zr => '0', ng => '0'),
        (x => "1001111011111000", y => "1000000011100001", zx => '1', nx => '0', zy => '1', ny => '1', f => '0', no => '0', o => "0000000000000000", zr => '1', ng => '0'),
        (x => "1101001110001110", y => "1111011111000111", zx => '1', nx => '0', zy => '0', ny => '0', f => '1', no => '0', o => "1111011111000111", zr => '0', ng => '1'),
        (x => "1100100100011110", y => "1010100010100100", zx => '1', nx => '1', zy => '1', ny => '1', f => '1', no => '1', o => "0000000000000001", zr => '0', ng => '0'),
        (x => "0111101000100000", y => "1011010100111101", zx => '1', nx => '0', zy => '1', ny => '0', f => '0', no => '1', o => "1111111111111111", zr => '0', ng => '1'),
        (x => "0110100101110010", y => "0101110110111000", zx => '0', nx => '0', zy => '0', ny => '0', f => '1', no => '1', o => "0011100011010101", zr => '0', ng => '0'),
        (x => "1101000101101001", y => "1001101110001000", zx => '1', nx => '0', zy => '0', ny => '0', f => '1', no => '1', o => "0110010001110111", zr => '0', ng => '0'),
        (x => "1101111010110000", y => "1100110110100101", zx => '0', nx => '1', zy => '1', ny => '0', f => '1', no => '0', o => "0010000101001111", zr => '0', ng => '0'),
        (x => "0110011100011000", y => "1001000000000101", zx => '0', nx => '0', zy => '1', ny => '0', f => '0', no => '1', o => "1111111111111111", zr => '0', ng => '1'),
        (x => "0110110111010100", y => "0111101110111011", zx => '0', nx => '0', zy => '1', ny => '1', f => '0', no => '0', o => "0110110111010100", zr => '0', ng => '0'),
        (x => "0000111111010011", y => "0111010100010010", zx => '0', nx => '1', zy => '1', ny => '1', f => '0', no => '0', o => "1111000000101100", zr => '0', ng => '1'),
        (x => "1011001001101101", y => "1010111110000111", zx => '0', nx => '1', zy => '1', ny => '1', f => '0', no => '0', o => "0100110110010010", zr => '0', ng => '0'),
        (x => "1100111001100001", y => "0101011011011111", zx => '1', nx => '0', zy => '1', ny => '0', f => '1', no => '1', o => "1111111111111111", zr => '0', ng => '1'),
        (x => "0110001100000010", y => "0111001010001001", zx => '0', nx => '1', zy => '0', ny => '0', f => '1', no => '1', o => "1111000001111001", zr => '0', ng => '1'),
        (x => "0010100011101100", y => "1011101000011100", zx => '1', nx => '0', zy => '1', ny => '1', f => '1', no => '1', o => "0000000000000000", zr => '1', ng => '0'),
        (x => "1010110000001000", y => "0001101001010110", zx => '0', nx => '1', zy => '0', ny => '1', f => '1', no => '0', o => "0011100110100000", zr => '0', ng => '0'),
        (x => "1100011011001101", y => "1001011000000100", zx => '0', nx => '0', zy => '1', ny => '0', f => '1', no => '1', o => "0011100100110010", zr => '0', ng => '0'),
        (x => "0000100110010100", y => "1111111111010111", zx => '0', nx => '1', zy => '1', ny => '0', f => '0', no => '1', o => "1111111111111111", zr => '0', ng => '1'),
        (x => "0011000111110000", y => "1111011100111101", zx => '0', nx => '1', zy => '0', ny => '0', f => '0', no => '1', o => "0011100111110010", zr => '0', ng => '0'),
        (x => "0010100011011000", y => "1110010111000101", zx => '0', nx => '0', zy => '0', ny => '1', f => '0', no => '0', o => "0000100000011000", zr => '0', ng => '0'),
        (x => "0001100100011010", y => "0001011010101001", zx => '0', nx => '1', zy => '0', ny => '1', f => '1', no => '0', o => "1101000000111011", zr => '0', ng => '1'),
        (x => "0100110010111001", y => "0000111101100000", zx => '0', nx => '1', zy => '0', ny => '0', f => '0', no => '0', o => "0000001101000000", zr => '0', ng => '0'),
        (x => "1000010111111101", y => "1000110110101111", zx => '1', nx => '0', zy => '0', ny => '0', f => '1', no => '0', o => "1000110110101111", zr => '0', ng => '1'),
        (x => "1001000111100011", y => "1100011010110000", zx => '0', nx => '0', zy => '1', ny => '0', f => '1', no => '0', o => "1001000111100011", zr => '0', ng => '1'),
        (x => "0000010111011100", y => "0100111001100011", zx => '1', nx => '1', zy => '0', ny => '1', f => '1', no => '1', o => "0100111001100100", zr => '0', ng => '0'),
        (x => "0111111101011000", y => "0001001010000111", zx => '1', nx => '1', zy => '1', ny => '1', f => '1', no => '1', o => "0000000000000001", zr => '0', ng => '0'),
        (x => "0101001100100000", y => "0100100110100111", zx => '0', nx => '0', zy => '0', ny => '1', f => '0', no => '1', o => "1110110111111111", zr => '0', ng => '1'),
        (x => "1000000100110001", y => "1111101011110001", zx => '1', nx => '1', zy => '0', ny => '1', f => '1', no => '0', o => "0000010100001101", zr => '0', ng => '0'),
        (x => "1100000110111100", y => "0010011100011100", zx => '0', nx => '1', zy => '1', ny => '1', f => '1', no => '0', o => "0011111001000010", zr => '0', ng => '0'),
        (x => "0010000011101110", y => "0010110101101001", zx => '1', nx => '0', zy => '0', ny => '1', f => '0', no => '0', o => "0000000000000000", zr => '1', ng => '0'),
        (x => "0010011001010000", y => "1000101001111010", zx => '1', nx => '1', zy => '1', ny => '0', f => '0', no => '1', o => "1111111111111111", zr => '0', ng => '1'),
        (x => "1110010010011001", y => "0001001011111111", zx => '1', nx => '1', zy => '1', ny => '0', f => '1', no => '1', o => "0000000000000000", zr => '1', ng => '0'),
        (x => "1110011000010110", y => "0110001001001110", zx => '0', nx => '1', zy => '1', ny => '0', f => '1', no => '1', o => "1110011000010110", zr => '0', ng => '1'),
        (x => "0001011110000000", y => "1011000010010010", zx => '1', nx => '1', zy => '0', ny => '1', f => '1', no => '1', o => "1011000010010011", zr => '0', ng => '1'),
        (x => "1100011111001110", y => "1000010110011110", zx => '0', nx => '1', zy => '0', ny => '0', f => '0', no => '1', o => "1111111111101111", zr => '0', ng => '1'),
        (x => "1000011001100000", y => "0110010000011000", zx => '1', nx => '1', zy => '0', ny => '1', f => '0', no => '0', o => "1001101111100111", zr => '0', ng => '1'),
        (x => "0100001110101011", y => "1111100111100110", zx => '1', nx => '0', zy => '1', ny => '0', f => '0', no => '0', o => "0000000000000000", zr => '1', ng => '0'),
        (x => "1100101001111111", y => "1001100111011101", zx => '1', nx => '0', zy => '1', ny => '1', f => '0', no => '0', o => "0000000000000000", zr => '1', ng => '0'),
        (x => "1101101111001000", y => "1101101011101001", zx => '1', nx => '0', zy => '1', ny => '0', f => '1', no => '0', o => "0000000000000000", zr => '1', ng => '0'),
        (x => "1110001011010100", y => "1100000110001100", zx => '1', nx => '0', zy => '1', ny => '0', f => '1', no => '1', o => "1111111111111111", zr => '0', ng => '1'),
        (x => "0011000000011001", y => "1001010101100011", zx => '0', nx => '0', zy => '0', ny => '0', f => '1', no => '0', o => "1100010101111100", zr => '0', ng => '1'),
        (x => "0111101011010101", y => "0001010101101001", zx => '0', nx => '1', zy => '1', ny => '0', f => '1', no => '0', o => "1000010100101010", zr => '0', ng => '1'),
        (x => "1011011110111010", y => "1001110011001100", zx => '0', nx => '0', zy => '0', ny => '0', f => '1', no => '0', o => "0101010010000110", zr => '0', ng => '0'),
        (x => "1111001011100100", y => "1011110000010011", zx => '0', nx => '0', zy => '1', ny => '0', f => '0', no => '1', o => "1111111111111111", zr => '0', ng => '1'),
        (x => "1010100010110101", y => "0001011101010110", zx => '0', nx => '0', zy => '0', ny => '1', f => '0', no => '1', o => "0101011101011110", zr => '0', ng => '0'),
        (x => "0101101101110001", y => "1010001101011111", zx => '1', nx => '1', zy => '1', ny => '1', f => '0', no => '1', o => "0000000000000000", zr => '1', ng => '0'),
        (x => "0101001011111010", y => "1010000011001001", zx => '1', nx => '1', zy => '1', ny => '0', f => '0', no => '0', o => "0000000000000000", zr => '1', ng => '0'),
        (x => "1101010010110010", y => "0111000100100011", zx => '0', nx => '0', zy => '1', ny => '0', f => '1', no => '0', o => "1101010010110010", zr => '0', ng => '1'),
        (x => "1110111010001010", y => "0001111111001100", zx => '1', nx => '1', zy => '0', ny => '1', f => '0', no => '1', o => "0001111111001100", zr => '0', ng => '0'),
        (x => "1111101001100101", y => "0001111100100111", zx => '0', nx => '1', zy => '0', ny => '1', f => '0', no => '1', o => "1111111101100111", zr => '0', ng => '1'),
        (x => "0011011101110010", y => "1111000001110010", zx => '0', nx => '0', zy => '1', ny => '1', f => '1', no => '0', o => "0011011101110001", zr => '0', ng => '0'),
        (x => "0111010011010110", y => "0010100101101100", zx => '0', nx => '1', zy => '0', ny => '0', f => '1', no => '1', o => "0100101101101010", zr => '0', ng => '0'),
        (x => "1010110111011110", y => "1010101110101001", zx => '1', nx => '1', zy => '0', ny => '0', f => '0', no => '1', o => "0101010001010110", zr => '0', ng => '0'),
        (x => "0100111100101000", y => "0101110101000001", zx => '0', nx => '1', zy => '0', ny => '1', f => '1', no => '0', o => "0101001110010101", zr => '0', ng => '0'),
        (x => "0001101010011111", y => "1110001110100000", zx => '0', nx => '0', zy => '1', ny => '0', f => '0', no => '1', o => "1111111111111111", zr => '0', ng => '1'),
        (x => "0010110011110110", y => "1010011000101110", zx => '1', nx => '1', zy => '1', ny => '0', f => '0', no => '1', o => "1111111111111111", zr => '0', ng => '1'),
        (x => "0010011110010111", y => "1111001011000101", zx => '0', nx => '0', zy => '1', ny => '0', f => '1', no => '0', o => "0010011110010111", zr => '0', ng => '0'),
        (x => "0010100000001001", y => "1001111100000110", zx => '1', nx => '1', zy => '0', ny => '1', f => '1', no => '0', o => "0110000011111000", zr => '0', ng => '0'),
        (x => "1100011011011010", y => "0111110001000010", zx => '0', nx => '1', zy => '1', ny => '0', f => '0', no => '0', o => "0000000000000000", zr => '1', ng => '0'),
        (x => "1010111100100011", y => "0101111111001110", zx => '0', nx => '1', zy => '0', ny => '1', f => '0', no => '0', o => "0000000000010000", zr => '0', ng => '0')
    );

    FUNCTION slv_to_string (slv : STD_LOGIC_VECTOR) RETURN STRING IS
        VARIABLE str : STRING (slv'length - 1 DOWNTO 1) := (OTHERS => NUL);
    BEGIN
        FOR n IN slv'length - 1 DOWNTO 1 LOOP
            str(n) := STD_LOGIC'image(slv((n - 1)))(2);
        END LOOP;
        RETURN str;
    END FUNCTION;

BEGIN
    bench : my_alu PORT MAP(x, y, zx, nx, zy, ny, f, no, o_actual, zr_actual, ng_actual);

    PROCESS
    BEGIN

        FOR n IN test_cases'RANGE LOOP
            x <= test_cases(n).x;
            y <= test_cases(n).y;
            zx <= test_cases(n).zx;
            nx <= test_cases(n).nx;
            zy <= test_cases(n).zy;
            ny <= test_cases(n).ny;
            f <= test_cases(n).f;
            no <= test_cases(n).no;
            o_expected <= test_cases(n).o;
            zr_expected <= test_cases(n).zr;
            ng_expected <= test_cases(n).ng;

            WAIT FOR 10 ns;

            ASSERT (o_actual = o_expected AND zr_actual = zr_expected AND ng_actual = ng_expected)
            REPORT "test failed for " &
                "x = " & slv_to_string(x) &
                ", y = " & slv_to_string(y) &
                ", zx = " & STD_LOGIC'image(zx) &
                ", nx = " & STD_LOGIC'image(nx) &
                ", zy = " & STD_LOGIC'image(zy) &
                ", ny = " & STD_LOGIC'image(ny) &
                ", f = " & STD_LOGIC'image(f) &
                ", no = " & STD_LOGIC'image(no) &
                ". expected o = " & slv_to_string(o_expected) &
                ", got " & slv_to_string(o_actual) &
                ". expected zr = " & STD_LOGIC'image(zr_expected) &
                ", got " & STD_LOGIC'image(zr_actual) &
                ". expected ng = " & STD_LOGIC'image(ng_expected) &
                ", got " & STD_LOGIC'image(ng_actual) SEVERITY error;
        END LOOP;
        WAIT;

    END PROCESS;

END behavioral;