LIBRARY ieee;
USE ieee.std_logic_1164.ALL;

ENTITY my_ram512_testbench IS
END my_ram512_testbench;

ARCHITECTURE behavioral OF my_ram512_testbench IS
    COMPONENT my_ram512
        PORT (
            clk : IN STD_LOGIC;
            load : IN STD_LOGIC;
            i : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
            sel : IN STD_LOGIC_VECTOR (8 DOWNTO 0);
            o : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
        );
    END COMPONENT;

    SIGNAL previous : STD_LOGIC_VECTOR (15 DOWNTO 0);
    SIGNAL clk : STD_LOGIC;
    SIGNAL load : STD_LOGIC;
    SIGNAL i : STD_LOGIC_VECTOR (15 DOWNTO 0);
    SIGNAL sel : STD_LOGIC_VECTOR (8 DOWNTO 0);
    SIGNAL o_actual : STD_LOGIC_VECTOR (15 DOWNTO 0);
    SIGNAL o_expected : STD_LOGIC_VECTOR (15 DOWNTO 0);

    CONSTANT clk_period : TIME := 10 ns;

    TYPE test_case IS RECORD
        previous : STD_LOGIC_VECTOR (15 DOWNTO 0);
        load : STD_LOGIC;
        i : STD_LOGIC_VECTOR (15 DOWNTO 0);
        sel : STD_LOGIC_VECTOR (8 DOWNTO 0);
        o : STD_LOGIC_VECTOR (15 DOWNTO 0);
    END RECORD;

    TYPE test_case_array IS ARRAY (NATURAL RANGE <>) OF test_case;
    CONSTANT test_cases : test_case_array := (
        -- previous, load, i, sel, o
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "1110001000000100", sel => "001101011", o => "UUUUUUUUUUUUUUUU"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "1100111000001100", sel => "010110011", o => "UUUUUUUUUUUUUUUU"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "1100011000100101", sel => "010100111", o => "UUUUUUUUUUUUUUUU"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "0011111111011011", sel => "010110100", o => "UUUUUUUUUUUUUUUU"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "0111010111101011", sel => "001100111", o => "UUUUUUUUUUUUUUUU"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "0001110111011101", sel => "011101000", o => "0001110111011101"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "0100100011011000", sel => "000101100", o => "0100100011011000"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "1011001000000000", sel => "011010101", o => "UUUUUUUUUUUUUUUU"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "0000000111001100", sel => "000011011", o => "UUUUUUUUUUUUUUUU"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "0101000111101111", sel => "010110001", o => "UUUUUUUUUUUUUUUU"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "1110110101011010", sel => "001111110", o => "1110110101011010"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "0111001100001110", sel => "001111010", o => "0111001100001110"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "0100011010110101", sel => "000101010", o => "UUUUUUUUUUUUUUUU"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "0101010101101001", sel => "000111011", o => "UUUUUUUUUUUUUUUU"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "1100110111010001", sel => "000101011", o => "1100110111010001"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "0111101110111001", sel => "000001101", o => "UUUUUUUUUUUUUUUU"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "0100001111100110", sel => "001111000", o => "UUUUUUUUUUUUUUUU"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "0100000110111011", sel => "010110001", o => "0100000110111011"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "0010010011010110", sel => "010110011", o => "0010010011010110"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "0010100110000111", sel => "010111110", o => "0010100110000111"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "0100010100000101", sel => "001011010", o => "0100010100000101"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "0001111110000000", sel => "011111011", o => "0001111110000000"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "0110010110101010", sel => "010101001", o => "0110010110101010"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "0110101011100101", sel => "001111011", o => "UUUUUUUUUUUUUUUU"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "1010111000010000", sel => "000101001", o => "1010111000010000"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "0001011100011101", sel => "011000010", o => "0001011100011101"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "0100101010010101", sel => "000111001", o => "0100101010010101"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "1111000001000110", sel => "010000111", o => "UUUUUUUUUUUUUUUU"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "1110101011111010", sel => "011010110", o => "UUUUUUUUUUUUUUUU"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "1000111010111000", sel => "011110010", o => "1000111010111000"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "0101111100010010", sel => "011111101", o => "UUUUUUUUUUUUUUUU"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "0011111000001110", sel => "001100010", o => "UUUUUUUUUUUUUUUU"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "1111100110110111", sel => "011010110", o => "1111100110110111"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "0101100000110010", sel => "011111111", o => "UUUUUUUUUUUUUUUU"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "1001100101011100", sel => "010010001", o => "1001100101011100"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "0011001100011110", sel => "011110101", o => "UUUUUUUUUUUUUUUU"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "0100001101010111", sel => "000010010", o => "UUUUUUUUUUUUUUUU"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "0001001011011111", sel => "000010101", o => "UUUUUUUUUUUUUUUU"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "0101001110110101", sel => "011010011", o => "UUUUUUUUUUUUUUUU"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "0000011110100111", sel => "001100111", o => "UUUUUUUUUUUUUUUU"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "1000000010100100", sel => "010000010", o => "1000000010100100"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "1010110000000111", sel => "010100010", o => "1010110000000111"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "1111110011011101", sel => "001000011", o => "UUUUUUUUUUUUUUUU"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "1011100111011100", sel => "010001110", o => "UUUUUUUUUUUUUUUU"),
        (previous => "0010100110000111", load => '0', i => "0011100001101101", sel => "010111110", o => "0010100110000111"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "0100011001100010", sel => "011111111", o => "0100011001100010"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "0101111101110100", sel => "001011110", o => "UUUUUUUUUUUUUUUU"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "1100011110001001", sel => "001010010", o => "1100011110001001"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "1100000001011100", sel => "010001100", o => "1100000001011100"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "0110111011000011", sel => "011000001", o => "UUUUUUUUUUUUUUUU"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "1111110001000101", sel => "010101101", o => "1111110001000101"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "1010110111101000", sel => "010101100", o => "UUUUUUUUUUUUUUUU"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "1010001100101011", sel => "010111001", o => "1010001100101011"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "0100000110111001", sel => "001111101", o => "0100000110111001"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "1111010001110111", sel => "001110100", o => "UUUUUUUUUUUUUUUU"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "0110100101110111", sel => "011000110", o => "0110100101110111"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "1011011111010101", sel => "000110111", o => "1011011111010101"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "0010101000100111", sel => "000000000", o => "0010101000100111"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "1011000010110011", sel => "010100111", o => "1011000010110011"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "0011011001110100", sel => "000000100", o => "0011011001110100"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "0100101000100010", sel => "000001001", o => "UUUUUUUUUUUUUUUU"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "0100101011001110", sel => "010110010", o => "UUUUUUUUUUUUUUUU"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "0111011010001000", sel => "001100010", o => "0111011010001000"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "1100011100000101", sel => "011101111", o => "UUUUUUUUUUUUUUUU"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "1001010001111001", sel => "001011000", o => "UUUUUUUUUUUUUUUU"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "0111100001000000", sel => "000101110", o => "0111100001000000"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "1010010101110111", sel => "001100111", o => "UUUUUUUUUUUUUUUU"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "0101111101110111", sel => "000010101", o => "0101111101110111"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "1011100100011111", sel => "001001100", o => "UUUUUUUUUUUUUUUU"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "0000011000100011", sel => "011011111", o => "0000011000100011"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "0100111000101100", sel => "000110110", o => "0100111000101100"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "0001000111011110", sel => "011010011", o => "0001000111011110"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "1111110101000000", sel => "001010111", o => "1111110101000000"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "0000110100101111", sel => "000000111", o => "0000110100101111"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "1111101110000111", sel => "001101111", o => "UUUUUUUUUUUUUUUU"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "0000000010110110", sel => "001001111", o => "UUUUUUUUUUUUUUUU"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "0110001100011101", sel => "010100110", o => "UUUUUUUUUUUUUUUU"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "1000001000110010", sel => "011010010", o => "1000001000110010"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "0010010101111110", sel => "000100101", o => "UUUUUUUUUUUUUUUU"),
        (previous => "0100100011011000", load => '0', i => "0000110101011110", sel => "000101100", o => "0100100011011000"),
        (previous => "1011000010110011", load => '0', i => "1010100010010100", sel => "010100111", o => "1011000010110011"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "1111001101100111", sel => "001000100", o => "1111001101100111"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "1001101110111111", sel => "010101111", o => "1001101110111111"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "0100010011000110", sel => "010100011", o => "0100010011000110"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "0011000000110101", sel => "010011100", o => "UUUUUUUUUUUUUUUU"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "0101001010000101", sel => "000001110", o => "UUUUUUUUUUUUUUUU"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "0001010100101011", sel => "011000001", o => "UUUUUUUUUUUUUUUU"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "0010111111111110", sel => "011101011", o => "UUUUUUUUUUUUUUUU"),
        (previous => "1100000001011100", load => '1', i => "1100110100100011", sel => "010001100", o => "1100110100100011"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "1001110101001111", sel => "001001101", o => "1001110101001111"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "1101011011110110", sel => "000110001", o => "1101011011110110"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "1100010000111010", sel => "001000001", o => "1100010000111010"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "1010111111101010", sel => "000110000", o => "UUUUUUUUUUUUUUUU"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "0001000010001101", sel => "001100000", o => "UUUUUUUUUUUUUUUU"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "1010110100101001", sel => "010111111", o => "1010110100101001"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "0001101000110111", sel => "010100101", o => "UUUUUUUUUUUUUUUU"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "1100111111111000", sel => "001000010", o => "UUUUUUUUUUUUUUUU"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "0111001111100011", sel => "011111100", o => "UUUUUUUUUUUUUUUU"),
        (previous => "0001110111011101", load => '1', i => "0110010101110000", sel => "011101000", o => "0110010101110000"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "0101110110111101", sel => "001010011", o => "0101110110111101"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "0110001011101110", sel => "000011100", o => "0110001011101110"),
        (previous => "0111001100001110", load => '0', i => "1100001100101111", sel => "001111010", o => "0111001100001110"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "1001000001100000", sel => "000111111", o => "UUUUUUUUUUUUUUUU"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "1100011111000000", sel => "011000011", o => "1100011111000000"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "0111011001111111", sel => "000001101", o => "UUUUUUUUUUUUUUUU"),
        (previous => "1100110100100011", load => '1', i => "1001100000100100", sel => "010001100", o => "1001100000100100"),
        (previous => "1001100101011100", load => '0', i => "0010110101100110", sel => "010010001", o => "1001100101011100"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "1001100101100010", sel => "011000001", o => "1001100101100010"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "0101111001001011", sel => "011101111", o => "0101111001001011"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "1010000110011110", sel => "001000000", o => "UUUUUUUUUUUUUUUU"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "0111000010111011", sel => "011100001", o => "UUUUUUUUUUUUUUUU"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "0111010000110101", sel => "001111001", o => "UUUUUUUUUUUUUUUU"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "1001111101110100", sel => "001001011", o => "UUUUUUUUUUUUUUUU"),
        (previous => "0000110100101111", load => '0', i => "1000111000110111", sel => "000000111", o => "0000110100101111"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "1000010101000100", sel => "001010000", o => "1000010101000100"),
        (previous => "0001011100011101", load => '1', i => "1011010011010000", sel => "011000010", o => "1011010011010000"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "0110111101100001", sel => "001101011", o => "UUUUUUUUUUUUUUUU"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "1100101000100010", sel => "000001101", o => "UUUUUUUUUUUUUUUU"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "1111010100010001", sel => "010010011", o => "1111010100010001"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "1011110101010010", sel => "010001000", o => "UUUUUUUUUUUUUUUU"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "1100000000110011", sel => "000111011", o => "1100000000110011"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "1101010010101100", sel => "011011011", o => "UUUUUUUUUUUUUUUU"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "1011111011110111", sel => "010101011", o => "UUUUUUUUUUUUUUUU"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "0010111011111110", sel => "011011011", o => "0010111011111110"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "0011010101001110", sel => "011001011", o => "0011010101001110"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "0111111100010000", sel => "000111010", o => "0111111100010000"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "0010011001111100", sel => "011001110", o => "0010011001111100"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "1111101110001001", sel => "011001000", o => "1111101110001001"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "0111001000011100", sel => "000100100", o => "0111001000011100"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "1110111110100101", sel => "011001100", o => "1110111110100101"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "1101000111100000", sel => "000010010", o => "UUUUUUUUUUUUUUUU"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "0111101110111011", sel => "000010011", o => "0111101110111011"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "1011000001100111", sel => "001001001", o => "UUUUUUUUUUUUUUUU"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "0000000001000010", sel => "011110011", o => "0000000001000010"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "0011001100001110", sel => "011010100", o => "0011001100001110"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "1011111101001000", sel => "011111001", o => "UUUUUUUUUUUUUUUU"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "0011110100010110", sel => "011101110", o => "UUUUUUUUUUUUUUUU"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "1101100111011110", sel => "001000101", o => "1101100111011110"),
        (previous => "1010110100101001", load => '0', i => "0010111100000011", sel => "010111111", o => "1010110100101001"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "1001101011001111", sel => "001001010", o => "1001101011001111"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "1011111011100001", sel => "000100111", o => "1011111011100001"),
        (previous => "1011011111010101", load => '0', i => "0000101111110100", sel => "000110111", o => "1011011111010101"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "1111011000111101", sel => "011110100", o => "1111011000111101"),
        (previous => "0110010110101010", load => '0', i => "0001110100110000", sel => "010101001", o => "0110010110101010"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "0000111100000100", sel => "001011100", o => "UUUUUUUUUUUUUUUU"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "0101000011111101", sel => "001011101", o => "UUUUUUUUUUUUUUUU"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "1001011111101011", sel => "001101111", o => "1001011111101011"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "0101001100110001", sel => "011111101", o => "0101001100110001"),
        (previous => "0101111101110111", load => '0', i => "0100110011110000", sel => "000010101", o => "0101111101110111"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "0111101000111010", sel => "001001001", o => "0111101000111010"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "1001100001100001", sel => "000100010", o => "UUUUUUUUUUUUUUUU"),
        (previous => "0010111011111110", load => '0', i => "0110011110011000", sel => "011011011", o => "0010111011111110"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "1011110010001101", sel => "001001111", o => "1011110010001101"),
        (previous => "1100110111010001", load => '1', i => "0101011000110110", sel => "000101011", o => "0101011000110110"),
        (previous => "0111101000111010", load => '1', i => "0110001110010010", sel => "001001001", o => "0110001110010010"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "0001100111101111", sel => "001110101", o => "UUUUUUUUUUUUUUUU"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "1111100001011111", sel => "011101001", o => "UUUUUUUUUUUUUUUU"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "0010010101011100", sel => "001110100", o => "0010010101011100"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "1001110001110001", sel => "011011110", o => "1001110001110001"),
        (previous => "1001101011001111", load => '1', i => "1100111110111010", sel => "001001010", o => "1100111110111010"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "1010111011011100", sel => "010000110", o => "UUUUUUUUUUUUUUUU"),
        (previous => "1010110000000111", load => '0', i => "0000101110110111", sel => "010100010", o => "1010110000000111"),
        (previous => "0010010011010110", load => '1', i => "0110001000000111", sel => "010110011", o => "0110001000000111"),
        (previous => "0010101000100111", load => '1', i => "0110001000110010", sel => "000000000", o => "0110001000110010"),
        (previous => "1110110101011010", load => '1', i => "0000110001111011", sel => "001111110", o => "0000110001111011"),
        (previous => "0100011001100010", load => '1', i => "1001001111110000", sel => "011111111", o => "1001001111110000"),
        (previous => "0000110001111011", load => '0', i => "1011011111011001", sel => "001111110", o => "0000110001111011"),
        (previous => "0110010101110000", load => '0', i => "1011010101001110", sel => "011101000", o => "0110010101110000"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "0110011000101100", sel => "010000011", o => "UUUUUUUUUUUUUUUU"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "1111100101110110", sel => "000001110", o => "UUUUUUUUUUUUUUUU"),
        (previous => "0001000111011110", load => '1', i => "0000100111111100", sel => "011010011", o => "0000100111111100"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "0101011010011111", sel => "011111001", o => "UUUUUUUUUUUUUUUU"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "1110101101010010", sel => "010110111", o => "1110101101010010"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "1011111001010010", sel => "000000011", o => "1011111001010010"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "1110110011010000", sel => "010000100", o => "UUUUUUUUUUUUUUUU"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "1000010111010000", sel => "010011000", o => "UUUUUUUUUUUUUUUU"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "1101101001001110", sel => "010011011", o => "UUUUUUUUUUUUUUUU"),
        (previous => "0101001100110001", load => '0', i => "1000001000110110", sel => "011111101", o => "0101001100110001"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "1101000010111001", sel => "010111011", o => "UUUUUUUUUUUUUUUU"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "0001001011000111", sel => "011101011", o => "UUUUUUUUUUUUUUUU"),
        (previous => "1111100110110111", load => '1', i => "1100001010011010", sel => "011010110", o => "1100001010011010"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "0111100010010011", sel => "010011101", o => "UUUUUUUUUUUUUUUU"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "1001110001001010", sel => "000011011", o => "UUUUUUUUUUUUUUUU"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "1110101001001101", sel => "010100001", o => "UUUUUUUUUUUUUUUU"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "1011100011010010", sel => "001011000", o => "1011100011010010"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "0110101101101010", sel => "010001011", o => "0110101101101010"),
        (previous => "1111110001000101", load => '1', i => "0001110000000101", sel => "010101101", o => "0001110000000101"),
        (previous => "0110010110101010", load => '1', i => "1100001100000010", sel => "010101001", o => "1100001100000010"),
        (previous => "0000000001000010", load => '0', i => "1000010110111101", sel => "011110011", o => "0000000001000010"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "0000000010101001", sel => "001101001", o => "0000000010101001"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "0000001101111111", sel => "001010110", o => "0000001101111111"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "0011110100011100", sel => "000111111", o => "UUUUUUUUUUUUUUUU"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "1011100100110111", sel => "011000111", o => "UUUUUUUUUUUUUUUU"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "1101100111011000", sel => "010100001", o => "UUUUUUUUUUUUUUUU"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "0000000100110001", sel => "011001101", o => "UUUUUUUUUUUUUUUU"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "0011101110111100", sel => "011001010", o => "UUUUUUUUUUUUUUUU"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "0001110101101001", sel => "010010111", o => "0001110101101001"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "0101111000010011", sel => "010110010", o => "0101111000010011"),
        (previous => "1011111001010010", load => '0', i => "1011001100000110", sel => "000000011", o => "1011111001010010"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "1000001001110000", sel => "000001101", o => "1000001001110000"),
        (previous => "1001110001110001", load => '0', i => "1100010111000110", sel => "011011110", o => "1001110001110001"),
        (previous => "0110001110010010", load => '0', i => "1000011100000101", sel => "001001001", o => "0110001110010010"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "0001110011001100", sel => "001000111", o => "UUUUUUUUUUUUUUUU"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "0111001001101101", sel => "010010000", o => "UUUUUUUUUUUUUUUU"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "0100011000111010", sel => "000100110", o => "0100011000111010"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "1000010100000101", sel => "010001110", o => "1000010100000101"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "1011010010011100", sel => "001100000", o => "1011010010011100"),
        (previous => "1011011111010101", load => '0', i => "1010111101001111", sel => "000110111", o => "1011011111010101"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "1111011101010010", sel => "000010000", o => "UUUUUUUUUUUUUUUU"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "0101110101100000", sel => "010100110", o => "UUUUUUUUUUUUUUUU"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "1111010000111110", sel => "011100110", o => "UUUUUUUUUUUUUUUU"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "0111111010001000", sel => "010100100", o => "0111111010001000"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "0111010011001111", sel => "001111111", o => "0111010011001111"),
        (previous => "1001100101011100", load => '0', i => "0111001101011111", sel => "010010001", o => "1001100101011100"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "0110010010000101", sel => "001111011", o => "0110010010000101"),
        (previous => "0001110101101001", load => '0', i => "0000000100010011", sel => "010010111", o => "0001110101101001"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "1011010001110011", sel => "001101110", o => "UUUUUUUUUUUUUUUU"),
        (previous => "1001101110111111", load => '1', i => "1001101010101010", sel => "010101111", o => "1001101010101010"),
        (previous => "1011111001010010", load => '0', i => "0111011010111010", sel => "000000011", o => "1011111001010010"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "1100111001100001", sel => "001011110", o => "UUUUUUUUUUUUUUUU"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "1010001001000111", sel => "000101000", o => "UUUUUUUUUUUUUUUU"),
        (previous => "1010001100101011", load => '0', i => "1111010111101011", sel => "010111001", o => "1010001100101011"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "0000011001101010", sel => "001001110", o => "UUUUUUUUUUUUUUUU"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "1000110011111011", sel => "010110000", o => "1000110011111011"),
        (previous => "0000110001111011", load => '1', i => "0110001101110111", sel => "001111110", o => "0110001101110111"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "1000101100001110", sel => "010000111", o => "UUUUUUUUUUUUUUUU"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "0011111101111100", sel => "010010101", o => "UUUUUUUUUUUUUUUU"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "1001111000101100", sel => "001000000", o => "UUUUUUUUUUUUUUUU"),
        (previous => "0100101010010101", load => '1', i => "0000010100101111", sel => "000111001", o => "0000010100101111"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "0010011110001101", sel => "010000101", o => "UUUUUUUUUUUUUUUU"),
        (previous => "1101011011110110", load => '1', i => "1000011110110110", sel => "000110001", o => "1000011110110110"),
        (previous => "0110001011101110", load => '0', i => "1110101101101111", sel => "000011100", o => "0110001011101110"),
        (previous => "1000010100000101", load => '1', i => "1101100110111101", sel => "010001110", o => "1101100110111101"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "0110111101101101", sel => "011010000", o => "UUUUUUUUUUUUUUUU"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "0001111011101100", sel => "001110010", o => "0001111011101100"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "0010111001110011", sel => "010011001", o => "0010111001110011"),
        (previous => "0000100111111100", load => '0', i => "0010001100001001", sel => "011010011", o => "0000100111111100"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "1011000101001001", sel => "010000001", o => "UUUUUUUUUUUUUUUU"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "1000100010000010", sel => "011011010", o => "1000100010000010"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "1010000000001000", sel => "011101101", o => "1010000000001000"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "0101010100111001", sel => "001100001", o => "0101010100111001"),
        (previous => "0110001011101110", load => '0', i => "1001110001010101", sel => "000011100", o => "0110001011101110"),
        (previous => "1011010011010000", load => '1', i => "1111001111100100", sel => "011000010", o => "1111001111100100"),
        (previous => "0000100111111100", load => '1', i => "1101000010110100", sel => "011010011", o => "1101000010110100"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "1010011000100110", sel => "011100000", o => "1010011000100110"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "1101100010111111", sel => "001100011", o => "UUUUUUUUUUUUUUUU"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "0110100110010011", sel => "011110101", o => "0110100110010011"),
        (previous => "1011111001010010", load => '0', i => "0000110100010100", sel => "000000011", o => "1011111001010010"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "0101110111101110", sel => "000111101", o => "0101110111101110"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "1101001011011011", sel => "010100110", o => "1101001011011011"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "0011101000111100", sel => "010011101", o => "UUUUUUUUUUUUUUUU"),
        (previous => "1100111110111010", load => '0', i => "0011011001011000", sel => "001001010", o => "1100111110111010"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "1011110100011011", sel => "001100110", o => "UUUUUUUUUUUUUUUU"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "1101010011101110", sel => "001000000", o => "UUUUUUUUUUUUUUUU"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "0000101011001110", sel => "010000111", o => "0000101011001110"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "1100001000110010", sel => "010111010", o => "UUUUUUUUUUUUUUUU"),
        (previous => "1011010010011100", load => '1', i => "1000011000100111", sel => "001100000", o => "1000011000100111"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "1001011000101010", sel => "000010000", o => "UUUUUUUUUUUUUUUU"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "1001000001100111", sel => "000001000", o => "UUUUUUUUUUUUUUUU"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "0111101000001101", sel => "010000011", o => "UUUUUUUUUUUUUUUU"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "0111101010101011", sel => "000000110", o => "UUUUUUUUUUUUUUUU"),
        (previous => "1100011111000000", load => '1', i => "0001100111110101", sel => "011000011", o => "0001100111110101"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "0100001101011100", sel => "011010101", o => "UUUUUUUUUUUUUUUU"),
        (previous => "0011010101001110", load => '0', i => "1101000010011100", sel => "011001011", o => "0011010101001110"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "0011000100100011", sel => "001110101", o => "0011000100100011"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "1000001111011101", sel => "001000110", o => "1000001111011101"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "1111011100111101", sel => "011010111", o => "UUUUUUUUUUUUUUUU"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "1010111001001101", sel => "011111010", o => "UUUUUUUUUUUUUUUU"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "0101101001010110", sel => "000110010", o => "0101101001010110"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "1000001111011001", sel => "001011001", o => "UUUUUUUUUUUUUUUU"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "1100101011100000", sel => "001011011", o => "1100101011100000"),
        (previous => "0010111001110011", load => '1', i => "1000010010100011", sel => "010011001", o => "1000010010100011"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "0100110101111000", sel => "000110000", o => "0100110101111000"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "0001100101000011", sel => "011100010", o => "0001100101000011"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "1011100010111000", sel => "010000011", o => "UUUUUUUUUUUUUUUU"),
        (previous => "1000111010111000", load => '1', i => "1101000111111111", sel => "011110010", o => "1101000111111111"),
        (previous => "1111010100010001", load => '0', i => "0011110111010110", sel => "010010011", o => "1111010100010001"),
        (previous => "1100101011100000", load => '0', i => "0110010111010000", sel => "001011011", o => "1100101011100000"),
        (previous => "1001110101001111", load => '0', i => "0101011100000011", sel => "001001101", o => "1001110101001111"),
        (previous => "1101001011011011", load => '1', i => "0110111101011100", sel => "010100110", o => "0110111101011100"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "1000000110110111", sel => "000001100", o => "1000000110110111"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "1100100001010000", sel => "000011110", o => "UUUUUUUUUUUUUUUU"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "0111100110000001", sel => "000100101", o => "UUUUUUUUUUUUUUUU"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "0101001001100011", sel => "010001000", o => "0101001001100011"),
        (previous => "0000101011001110", load => '0', i => "0010011111100110", sel => "010000111", o => "0000101011001110"),
        (previous => "1100001100000010", load => '1', i => "0000010011011000", sel => "010101001", o => "0000010011011000"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "1010101101101011", sel => "010101000", o => "1010101101101011"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "1010000111000110", sel => "011100100", o => "1010000111000110"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "0111111000010011", sel => "001101110", o => "UUUUUUUUUUUUUUUU"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "1101000010111001", sel => "001001110", o => "UUUUUUUUUUUUUUUU"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "0001001111000110", sel => "000001000", o => "0001001111000110"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "1100000111100100", sel => "010100001", o => "UUUUUUUUUUUUUUUU"),
        (previous => "1001110001110001", load => '1', i => "1111010100001001", sel => "011011110", o => "1111010100001001"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "1111000010010001", sel => "010010010", o => "UUUUUUUUUUUUUUUU"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "1000010100011000", sel => "010001010", o => "1000010100011000"),
        (previous => "0111111100010000", load => '1', i => "1110001111000001", sel => "000111010", o => "1110001111000001"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "1001000001101001", sel => "011101001", o => "1001000001101001"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "1000001001001101", sel => "001101110", o => "1000001001001101"),
        (previous => "0001100111110101", load => '1', i => "0110011110111100", sel => "011000011", o => "0110011110111100"),
        (previous => "0110001011101110", load => '0', i => "1001101100001010", sel => "000011100", o => "0110001011101110"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "1010000000010010", sel => "011010000", o => "UUUUUUUUUUUUUUUU"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "0100000110110100", sel => "000111100", o => "UUUUUUUUUUUUUUUU"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "0000010010010010", sel => "011111000", o => "0000010010010010"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "0011011000100100", sel => "000110101", o => "UUUUUUUUUUUUUUUU"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "1110111110101110", sel => "011010101", o => "UUUUUUUUUUUUUUUU"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "1110100111101000", sel => "001011100", o => "1110100111101000"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "1111011011010001", sel => "010111100", o => "UUUUUUUUUUUUUUUU"),
        (previous => "0000101011001110", load => '0', i => "0101010000111111", sel => "010000111", o => "0000101011001110"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "0110100000000011", sel => "000011000", o => "UUUUUUUUUUUUUUUU"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "1000100100011111", sel => "010111101", o => "UUUUUUUUUUUUUUUU"),
        (previous => "0110001011101110", load => '1', i => "0010011011101111", sel => "000011100", o => "0010011011101111"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "1100001100101011", sel => "001000000", o => "1100001100101011"),
        (previous => "0110001110010010", load => '1', i => "0010011000100011", sel => "001001001", o => "0010011000100011"),
        (previous => "0100010100000101", load => '1', i => "1100100101011000", sel => "001011010", o => "1100100101011000"),
        (previous => "0101001100110001", load => '0', i => "1111111100101110", sel => "011111101", o => "0101001100110001"),
        (previous => "1110101101010010", load => '0', i => "1110111110001010", sel => "010110111", o => "1110101101010010"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "1001111101000110", sel => "000110011", o => "UUUUUUUUUUUUUUUU"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "1011100111001101", sel => "000010111", o => "1011100111001101"),
        (previous => "0010011000100011", load => '0', i => "1110000011100110", sel => "001001001", o => "0010011000100011"),
        (previous => "1011011111010101", load => '1', i => "1001001010100011", sel => "000110111", o => "1001001010100011"),
        (previous => "0100110101111000", load => '1', i => "1001111110111111", sel => "000110000", o => "1001111110111111"),
        (previous => "1100000000110011", load => '0', i => "0001110000000000", sel => "000111011", o => "1100000000110011"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "1100100101001001", sel => "011111010", o => "UUUUUUUUUUUUUUUU"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "1001110010100011", sel => "001001011", o => "UUUUUUUUUUUUUUUU"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "1000011010100000", sel => "011000000", o => "UUUUUUUUUUUUUUUU"),
        (previous => "1010000111000110", load => '1', i => "0000110001011000", sel => "011100100", o => "0000110001011000"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "0001000110001011", sel => "011110001", o => "0001000110001011"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "0010011010100010", sel => "011001111", o => "0010011010100010"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "1100110111101100", sel => "011101100", o => "1100110111101100"),
        (previous => "1000001001110000", load => '0', i => "0110111100100011", sel => "000001101", o => "1000001001110000"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "1010010101010011", sel => "001001100", o => "UUUUUUUUUUUUUUUU"),
        (previous => "0110010010000101", load => '0', i => "0001000010001110", sel => "001111011", o => "0110010010000101"),
        (previous => "1100001010011010", load => '1', i => "1111001010001000", sel => "011010110", o => "1111001010001000"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "0100111111010011", sel => "001010100", o => "UUUUUUUUUUUUUUUU"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "0101111010010100", sel => "000101010", o => "0101111010010100"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "0000111001111000", sel => "000101111", o => "0000111001111000"),
        (previous => "0010100110000111", load => '0', i => "0100100101101001", sel => "010111110", o => "0010100110000111"),
        (previous => "1111010100010001", load => '0', i => "0000011000111000", sel => "010010011", o => "1111010100010001"),
        (previous => "0100111000101100", load => '0', i => "1001100100100101", sel => "000110110", o => "0100111000101100"),
        (previous => "1010110100101001", load => '0', i => "0110101000110010", sel => "010111111", o => "1010110100101001"),
        (previous => "1100110111101100", load => '1', i => "0000001001111110", sel => "011101100", o => "0000001001111110"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "1000100011111010", sel => "011011000", o => "UUUUUUUUUUUUUUUU"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "1100000011010000", sel => "011000100", o => "UUUUUUUUUUUUUUUU"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "1101000000100100", sel => "011111001", o => "UUUUUUUUUUUUUUUU"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "1000000001001110", sel => "011010001", o => "UUUUUUUUUUUUUUUU"),
        (previous => "1100111110111010", load => '0', i => "1101000001111101", sel => "001001010", o => "1100111110111010"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "1011000000111011", sel => "000011011", o => "UUUUUUUUUUUUUUUU"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "1011111011001111", sel => "001110111", o => "UUUUUUUUUUUUUUUU"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "1011011000000101", sel => "001110110", o => "1011011000000101"),
        (previous => "1000011000100111", load => '1', i => "0111011011000101", sel => "001100000", o => "0111011011000101"),
        (previous => "1000001001001101", load => '0', i => "1001001110110001", sel => "001101110", o => "1000001001001101"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "1010110010001001", sel => "011010000", o => "UUUUUUUUUUUUUUUU"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "1101110101001101", sel => "011000000", o => "UUUUUUUUUUUUUUUU"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "1110111101000110", sel => "000111000", o => "UUUUUUUUUUUUUUUU"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "0111111100010111", sel => "010000100", o => "UUUUUUUUUUUUUUUU"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "0001001101100010", sel => "001100100", o => "UUUUUUUUUUUUUUUU"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "1011100001111101", sel => "010111101", o => "1011100001111101"),
        (previous => "0111010011001111", load => '0', i => "0111111111110101", sel => "001111111", o => "0111010011001111"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "1001000001101011", sel => "001111001", o => "UUUUUUUUUUUUUUUU"),
        (previous => "1000010010100011", load => '1', i => "1011011111001011", sel => "010011001", o => "1011011111001011"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "0110010100111010", sel => "011101010", o => "UUUUUUUUUUUUUUUU"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "0011111000001010", sel => "010111010", o => "0011111000001010"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "0101001011001010", sel => "010000100", o => "UUUUUUUUUUUUUUUU"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "1001011000000010", sel => "000011110", o => "UUUUUUUUUUUUUUUU"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "0101011110000111", sel => "011011100", o => "0101011110000111"),
        (previous => "1001000001101001", load => '1', i => "1111010111101011", sel => "011101001", o => "1111010111101011"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "0111111110101000", sel => "001110011", o => "0111111110101000"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "0011111000100111", sel => "000111000", o => "UUUUUUUUUUUUUUUU"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "0011011110100001", sel => "011001101", o => "0011011110100001"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "0000010100111010", sel => "001100111", o => "UUUUUUUUUUUUUUUU"),
        (previous => "0110100101110111", load => '0', i => "0001000100100100", sel => "011000110", o => "0110100101110111"),
        (previous => "1111001010001000", load => '0', i => "0101110111011111", sel => "011010110", o => "1111001010001000"),
        (previous => "1001011111101011", load => '0', i => "0111010001100011", sel => "001101111", o => "1001011111101011"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "0001010110000010", sel => "001010101", o => "0001010110000010"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "0001000101011110", sel => "010000001", o => "UUUUUUUUUUUUUUUU"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "1110100001000111", sel => "011000100", o => "1110100001000111"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "0110101010111010", sel => "001101010", o => "UUUUUUUUUUUUUUUU"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "0100100011110011", sel => "010001101", o => "0100100011110011"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "0100000111000000", sel => "010100101", o => "UUUUUUUUUUUUUUUU"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "0000101100100111", sel => "000101000", o => "UUUUUUUUUUUUUUUU"),
        (previous => "1011011000000101", load => '1', i => "0001101111101101", sel => "001110110", o => "0001101111101101"),
        (previous => "1001001111110000", load => '0', i => "0000011111000011", sel => "011111111", o => "1001001111110000"),
        (previous => "1001100101011100", load => '1', i => "0111101100110010", sel => "010010001", o => "0111101100110010"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "0101001110000111", sel => "011101110", o => "0101001110000111"),
        (previous => "1001110101001111", load => '0', i => "1000000000001000", sel => "001001101", o => "1001110101001111"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "0111111111001100", sel => "000110011", o => "0111111111001100"),
        (previous => "0011011001110100", load => '0', i => "0110011000110110", sel => "000000100", o => "0011011001110100"),
        (previous => "0110001101110111", load => '1', i => "1110101111000011", sel => "001111110", o => "1110101111000011"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "1001000001101000", sel => "000100000", o => "1001000001101000"),
        (previous => "0111011010001000", load => '0', i => "1110010010010000", sel => "001100010", o => "0111011010001000"),
        (previous => "0000011000100011", load => '1', i => "1010000000000111", sel => "011011111", o => "1010000000000111"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "0010100000000110", sel => "010000000", o => "UUUUUUUUUUUUUUUU"),
        (previous => "0110001000110010", load => '0', i => "1011101010010111", sel => "000000000", o => "0110001000110010"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "1010101010000101", sel => "011100011", o => "1010101010000101"),
        (previous => "0010011000100011", load => '1', i => "1000110111010010", sel => "001001001", o => "1000110111010010"),
        (previous => "1000001001110000", load => '1', i => "1011110000000101", sel => "000001101", o => "1011110000000101"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "0010101100001010", sel => "000011000", o => "UUUUUUUUUUUUUUUU"),
        (previous => "1111010100001001", load => '1', i => "0101101010001000", sel => "011011110", o => "0101101010001000"),
        (previous => "0001110101101001", load => '0', i => "1000100010101000", sel => "010010111", o => "0001110101101001"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "1110110100001011", sel => "000010000", o => "UUUUUUUUUUUUUUUU"),
        (previous => "1000110011111011", load => '1', i => "1000110011101010", sel => "010110000", o => "1000110011101010"),
        (previous => "0101110111101110", load => '1', i => "0111100101101010", sel => "000111101", o => "0111100101101010"),
        (previous => "0100100011110011", load => '1', i => "0001000001101010", sel => "010001101", o => "0001000001101010"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "1100011001001101", sel => "000001111", o => "UUUUUUUUUUUUUUUU"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "1011000010010110", sel => "000011000", o => "1011000010010110"),
        (previous => "1010111000010000", load => '0', i => "1110000010100011", sel => "000101001", o => "1010111000010000"),
        (previous => "0000110100101111", load => '0', i => "0011111010111100", sel => "000000111", o => "0000110100101111"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "0011010110011010", sel => "000011011", o => "0011010110011010"),
        (previous => "1101000111111111", load => '1', i => "0000111000110010", sel => "011110010", o => "0000111000110010"),
        (previous => "0101101001010110", load => '0', i => "0000101001000010", sel => "000110010", o => "0101101001010110"),
        (previous => "1011111001010010", load => '0', i => "0011010011110011", sel => "000000011", o => "1011111001010010"),
        (previous => "1000100010000010", load => '0', i => "1010101000110000", sel => "011011010", o => "1000100010000010"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "0111000110111110", sel => "010111000", o => "UUUUUUUUUUUUUUUU"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "0000011011001101", sel => "000101101", o => "UUUUUUUUUUUUUUUU"),
        (previous => "1011111011100001", load => '0', i => "1011110011100110", sel => "000100111", o => "1011111011100001"),
        (previous => "1111011000111101", load => '0', i => "0001010000001111", sel => "011110100", o => "1111011000111101"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "1000110000010110", sel => "011000111", o => "UUUUUUUUUUUUUUUU"),
        (previous => "0100010011000110", load => '0', i => "1000101100110001", sel => "010100011", o => "0100010011000110"),
        (previous => "0001001111000110", load => '0', i => "1111110100100100", sel => "000001000", o => "0001001111000110"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "0111001001010110", sel => "000010110", o => "0111001001010110"),
        (previous => "0111100001000000", load => '0', i => "1100111101011001", sel => "000101110", o => "0111100001000000"),
        (previous => "1000011110110110", load => '0', i => "1011010000110100", sel => "000110001", o => "1000011110110110"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "0100100011101100", sel => "010011101", o => "UUUUUUUUUUUUUUUU"),
        (previous => "0010010101011100", load => '0', i => "0100100000011001", sel => "001110100", o => "0010010101011100"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "0101110001000000", sel => "010011000", o => "UUUUUUUUUUUUUUUU"),
        (previous => "1100011110001001", load => '1', i => "0001001100110101", sel => "001010010", o => "0001001100110101"),
        (previous => "1000110011101010", load => '0', i => "0010100011111100", sel => "010110000", o => "1000110011101010"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "1100100010011111", sel => "011001010", o => "1100100010011111"),
        (previous => "0111010011001111", load => '1', i => "0100110010101000", sel => "001111111", o => "0100110010101000"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "0011110110111110", sel => "001100101", o => "UUUUUUUUUUUUUUUU"),
        (previous => "1101100110111101", load => '1', i => "1000100011101100", sel => "010001110", o => "1000100011101100"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "1011101100011101", sel => "010101010", o => "1011101100011101"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "0100110110111011", sel => "011110111", o => "0100110110111011"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "0101000100101111", sel => "000000001", o => "UUUUUUUUUUUUUUUU"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "1000101111000111", sel => "011011001", o => "1000101111000111"),
        (previous => "0001110101101001", load => '0', i => "1010111000011001", sel => "010010111", o => "0001110101101001"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "1001100011001010", sel => "001100101", o => "UUUUUUUUUUUUUUUU"),
        (previous => "1000110111010010", load => '1', i => "1000101010010100", sel => "001001001", o => "1000101010010100"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "1011100100010011", sel => "001011110", o => "1011100100010011"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "0011001001111001", sel => "010011000", o => "0011001001111001"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "0000000100000111", sel => "000101000", o => "UUUUUUUUUUUUUUUU"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "0101100110110010", sel => "000010001", o => "0101100110110010"),
        (previous => "0000111001111000", load => '0', i => "1110011010101001", sel => "000101111", o => "0000111001111000"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "0001100110101010", sel => "000111000", o => "0001100110101010"),
        (previous => "1100101011100000", load => '0', i => "1111100110000100", sel => "001011011", o => "1100101011100000"),
        (previous => "0010100110000111", load => '0', i => "0100001100011011", sel => "010111110", o => "0010100110000111"),
        (previous => "0000001101111111", load => '0', i => "0000101010000000", sel => "001010110", o => "0000001101111111"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "1101101111001001", sel => "011101010", o => "UUUUUUUUUUUUUUUU"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "0100001000101000", sel => "000011101", o => "UUUUUUUUUUUUUUUU"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "0011101011000000", sel => "011111001", o => "0011101011000000"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "0011011111101000", sel => "010010010", o => "UUUUUUUUUUUUUUUU"),
        (previous => "1011000010010110", load => '0', i => "0000100011111001", sel => "000011000", o => "1011000010010110"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "0110001000101000", sel => "010111100", o => "0110001000101000"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "1000110001100001", sel => "000011010", o => "UUUUUUUUUUUUUUUU"),
        (previous => "1010101101101011", load => '0', i => "1100111110111100", sel => "010101000", o => "1010101101101011"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "1000100001111010", sel => "011111100", o => "1000100001111010"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "1100100111010000", sel => "001101010", o => "UUUUUUUUUUUUUUUU"),
        (previous => "1010110000000111", load => '1', i => "1011110010111010", sel => "010100010", o => "1011110010111010"),
        (previous => "1001011111101011", load => '1', i => "0010100111010111", sel => "001101111", o => "0010100111010111"),
        (previous => "1011110010001101", load => '1', i => "0101110111010000", sel => "001001111", o => "0101110111010000"),
        (previous => "1010101101101011", load => '1', i => "1001011001100011", sel => "010101000", o => "1001011001100011"),
        (previous => "0001001111000110", load => '1', i => "0101110001111011", sel => "000001000", o => "0101110001111011"),
        (previous => "0011010110011010", load => '1', i => "0110101100110111", sel => "000011011", o => "0110101100110111"),
        (previous => "1111001010001000", load => '0', i => "0001000001010010", sel => "011010110", o => "1111001010001000"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "1001110011111010", sel => "000111100", o => "UUUUUUUUUUUUUUUU"),
        (previous => "0100011000111010", load => '0', i => "1001110011110110", sel => "000100110", o => "0100011000111010"),
        (previous => "0100100011011000", load => '0', i => "1011111001100001", sel => "000101100", o => "0100100011011000"),
        (previous => "0101111000010011", load => '0', i => "1001101000000011", sel => "010110010", o => "0101111000010011"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "1011101001110010", sel => "000000001", o => "UUUUUUUUUUUUUUUU"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "1101100011000001", sel => "001111001", o => "UUUUUUUUUUUUUUUU"),
        (previous => "1000110011101010", load => '1', i => "0010011101101001", sel => "010110000", o => "0010011101101001"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "1010011101110010", sel => "011010000", o => "1010011101110010"),
        (previous => "1111010111101011", load => '0', i => "1011001010001101", sel => "011101001", o => "1111010111101011"),
        (previous => "0101111010010100", load => '0', i => "0010111101100011", sel => "000101010", o => "0101111010010100"),
        (previous => "0011011110100001", load => '0', i => "0011011110100000", sel => "011001101", o => "0011011110100001"),
        (previous => "0101011000110110", load => '1', i => "1100010011000110", sel => "000101011", o => "1100010011000110"),
        (previous => "0011011001110100", load => '0', i => "0001100111110010", sel => "000000100", o => "0011011001110100"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "0100000110100100", sel => "010101100", o => "0100000110100100"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "0001011110100110", sel => "000001111", o => "UUUUUUUUUUUUUUUU"),
        (previous => "1000101010010100", load => '1', i => "1101111000011111", sel => "001001001", o => "1101111000011111"),
        (previous => "0101110110111101", load => '1', i => "1100111111001111", sel => "001010011", o => "1100111111001111"),
        (previous => "1001100101100010", load => '1', i => "0010010010011111", sel => "011000001", o => "0010010010011111"),
        (previous => "1011101100011101", load => '0', i => "1110010110001000", sel => "010101010", o => "1011101100011101"),
        (previous => "1100100010011111", load => '1', i => "0111010010110011", sel => "011001010", o => "0111010010110011"),
        (previous => "0111100101101010", load => '1', i => "0101111010000000", sel => "000111101", o => "0101111010000000"),
        (previous => "0000010011011000", load => '0', i => "0111001010101011", sel => "010101001", o => "0000010011011000"),
        (previous => "1000000110110111", load => '0', i => "0011100110101111", sel => "000001100", o => "1000000110110111"),
        (previous => "1010011101110010", load => '1', i => "0111110101011100", sel => "011010000", o => "0111110101011100"),
        (previous => "0011001001111001", load => '1', i => "1111101001101011", sel => "010011000", o => "1111101001101011"),
        (previous => "1000001000110010", load => '0', i => "1101101010110100", sel => "011010010", o => "1000001000110010"),
        (previous => "0011011110100001", load => '1', i => "0111110000000111", sel => "011001101", o => "0111110000000111"),
        (previous => "0101101001010110", load => '1', i => "0111010011001000", sel => "000110010", o => "0111010011001000"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "0010000101110010", sel => "000001001", o => "0010000101110010"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "1110110100111101", sel => "001101101", o => "UUUUUUUUUUUUUUUU"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "1110100001111010", sel => "000110101", o => "UUUUUUUUUUUUUUUU"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "1011000000100011", sel => "010011100", o => "UUUUUUUUUUUUUUUU"),
        (previous => "0111010010110011", load => '1', i => "1110000100110000", sel => "011001010", o => "1110000100110000"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "0011101000000000", sel => "011101011", o => "0011101000000000"),
        (previous => "0010011101101001", load => '0', i => "0101010010011000", sel => "010110000", o => "0010011101101001"),
        (previous => "0110101100110111", load => '0', i => "1110101101101010", sel => "000011011", o => "0110101100110111"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "1101011100111000", sel => "010100101", o => "UUUUUUUUUUUUUUUU"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "0011111101101010", sel => "011111110", o => "UUUUUUUUUUUUUUUU"),
        (previous => "0100110110111011", load => '1', i => "1100101101110100", sel => "011110111", o => "1100101101110100"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "0010110111100001", sel => "001111001", o => "UUUUUUUUUUUUUUUU"),
        (previous => "0001110000000101", load => '0', i => "1001011000010110", sel => "010101101", o => "0001110000000101"),
        (previous => "0111011010001000", load => '1', i => "0011101110110011", sel => "001100010", o => "0011101110110011"),
        (previous => "1111001111100100", load => '1', i => "1110001101111101", sel => "011000010", o => "1110001101111101"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "1010011101101000", sel => "011010001", o => "UUUUUUUUUUUUUUUU"),
        (previous => "0101111010000000", load => '0', i => "1100100100011000", sel => "000111101", o => "0101111010000000"),
        (previous => "0111101110111011", load => '1', i => "0110000000110011", sel => "000010011", o => "0110000000110011"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "0100101011011000", sel => "010011110", o => "0100101011011000"),
        (previous => "1001111110111111", load => '1', i => "0101100011010111", sel => "000110000", o => "0101100011010111"),
        (previous => "1000010100011000", load => '1', i => "1010111011001110", sel => "010001010", o => "1010111011001110"),
        (previous => "1111110101000000", load => '1', i => "0011001001000111", sel => "001010111", o => "0011001001000111"),
        (previous => "0101010100111001", load => '1', i => "0101011111110101", sel => "001100001", o => "0101011111110101"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "0111111001010111", sel => "011100101", o => "UUUUUUUUUUUUUUUU"),
        (previous => "0001000001101010", load => '0', i => "0001100000011001", sel => "010001101", o => "0001000001101010"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "0101111011101010", sel => "001100100", o => "UUUUUUUUUUUUUUUU"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "1101000000100111", sel => "000111100", o => "1101000000100111"),
        (previous => "0001110000000101", load => '0', i => "0110011000111011", sel => "010101101", o => "0001110000000101"),
        (previous => "0101001001100011", load => '1', i => "1111101111011001", sel => "010001000", o => "1111101111011001"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "0000110100001001", sel => "010011011", o => "UUUUUUUUUUUUUUUU"),
        (previous => "1011000010010110", load => '0', i => "0000111010010011", sel => "000011000", o => "1011000010010110"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "0010000111101011", sel => "000001010", o => "UUUUUUUUUUUUUUUU"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "0011010001001100", sel => "011011101", o => "0011010001001100"),
        (previous => "0110100101110111", load => '0', i => "0010111000110010", sel => "011000110", o => "0110100101110111"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "1011111110111111", sel => "001100011", o => "1011111110111111"),
        (previous => "0100000110111001", load => '1', i => "1100101000100011", sel => "001111101", o => "1100101000100011"),
        (previous => "1001001111110000", load => '1', i => "1000011101100000", sel => "011111111", o => "1000011101100000"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "0100110000001101", sel => "010011010", o => "UUUUUUUUUUUUUUUU"),
        (previous => "0000000010101001", load => '1', i => "0000001110010101", sel => "001101001", o => "0000001110010101"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "1000010100110000", sel => "000010000", o => "UUUUUUUUUUUUUUUU"),
        (previous => "1000100011101100", load => '1', i => "0001000001001000", sel => "010001110", o => "0001000001001000"),
        (previous => "1000100010000010", load => '0', i => "0111000001010010", sel => "011011010", o => "1000100010000010"),
        (previous => "1000001001001101", load => '1', i => "1101001100101111", sel => "001101110", o => "1101001100101111"),
        (previous => "1100101101110100", load => '1', i => "1100111011110110", sel => "011110111", o => "1100111011110110"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "1001111101011001", sel => "011010111", o => "UUUUUUUUUUUUUUUU"),
        (previous => "0111110101011100", load => '1', i => "0010011111010110", sel => "011010000", o => "0010011111010110"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "0000111111010101", sel => "010110100", o => "0000111111010101"),
        (previous => "1010110100101001", load => '0', i => "0010000001110000", sel => "010111111", o => "1010110100101001"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "1011100111011001", sel => "000000101", o => "1011100111011001"),
        (previous => "0111001000011100", load => '1', i => "0010011011101001", sel => "000100100", o => "0010011011101001"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "1100000001110111", sel => "001001100", o => "UUUUUUUUUUUUUUUU"),
        (previous => "0000110100101111", load => '0', i => "0011010101010001", sel => "000000111", o => "0000110100101111"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "1011011111000000", sel => "010101110", o => "UUUUUUUUUUUUUUUU"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "1001111110110111", sel => "010100001", o => "UUUUUUUUUUUUUUUU"),
        (previous => "0110100101110111", load => '1', i => "0110101110001111", sel => "011000110", o => "0110101110001111"),
        (previous => "1011101100011101", load => '1', i => "0011001101011111", sel => "010101010", o => "0011001101011111"),
        (previous => "0100000110111011", load => '0', i => "0101011000010011", sel => "010110001", o => "0100000110111011"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "1010001111010010", sel => "000011001", o => "UUUUUUUUUUUUUUUU"),
        (previous => "0001000001101010", load => '1', i => "1000001011010111", sel => "010001101", o => "1000001011010111"),
        (previous => "0001110101101001", load => '0', i => "1110111011111011", sel => "010010111", o => "0001110101101001"),
        (previous => "0010011111010110", load => '1', i => "1111010101000111", sel => "011010000", o => "1111010101000111"),
        (previous => "0001001100110101", load => '1', i => "1010010001001111", sel => "001010010", o => "1010010001001111"),
        (previous => "1011111011100001", load => '1', i => "0001110111111101", sel => "000100111", o => "0001110111111101"),
        (previous => "1100010011000110", load => '0', i => "1001011010011110", sel => "000101011", o => "1100010011000110"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "0011110001100100", sel => "000100101", o => "0011110001100100"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "1100111100001110", sel => "001111000", o => "1100111100001110"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "0001100010111111", sel => "010100001", o => "UUUUUUUUUUUUUUUU"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "1010000011011000", sel => "010011111", o => "1010000011011000"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "1011001101100110", sel => "000001110", o => "UUUUUUUUUUUUUUUU"),
        (previous => "0001010110000010", load => '0', i => "0101001111111101", sel => "001010101", o => "0001010110000010"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "0000011111001101", sel => "010000110", o => "0000011111001101"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "1101111100100000", sel => "000101101", o => "UUUUUUUUUUUUUUUU"),
        (previous => "0100011000111010", load => '1', i => "0100101001000111", sel => "000100110", o => "0100101001000111"),
        (previous => "1010000000000111", load => '1', i => "0001110001110010", sel => "011011111", o => "0001110001110010"),
        (previous => "1000010101000100", load => '1', i => "0010010010010111", sel => "001010000", o => "0010010010010111"),
        (previous => "0101110111010000", load => '1', i => "0000001000001111", sel => "001001111", o => "0000001000001111"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "1101110010110000", sel => "010101110", o => "1101110010110000"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "1100010001001111", sel => "000100001", o => "1100010001001111"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "1101100101011101", sel => "001100110", o => "1101100101011101"),
        (previous => "1000000010100100", load => '0', i => "1101010110110011", sel => "010000010", o => "1000000010100100"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "1110000000111001", sel => "010011010", o => "UUUUUUUUUUUUUUUU"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "1011100101100110", sel => "011111010", o => "UUUUUUUUUUUUUUUU"),
        (previous => "1001011001100011", load => '1', i => "1001011010001101", sel => "010101000", o => "1001011010001101"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "0010111101101100", sel => "001010100", o => "0010111101101100"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "0010001110111100", sel => "010011101", o => "UUUUUUUUUUUUUUUU"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "1101111100001100", sel => "001001011", o => "1101111100001100"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "1001010010111010", sel => "000000110", o => "1001010010111010"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "1001101011011011", sel => "010000001", o => "UUUUUUUUUUUUUUUU"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "1001010101000001", sel => "011010101", o => "UUUUUUUUUUUUUUUU"),
        (previous => "0001000001001000", load => '1', i => "0000011011000100", sel => "010001110", o => "0000011011000100"),
        (previous => "1101100111011110", load => '0', i => "1101111001011110", sel => "001000101", o => "1101100111011110"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "0001000101011000", sel => "011001001", o => "UUUUUUUUUUUUUUUU"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "0100010000000001", sel => "001101101", o => "0100010000000001"),
        (previous => "1011100011010010", load => '0', i => "1001010001010101", sel => "001011000", o => "1011100011010010"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "1001100011110010", sel => "010110101", o => "UUUUUUUUUUUUUUUU"),
        (previous => "0000010011011000", load => '0', i => "1000111000111101", sel => "010101001", o => "0000010011011000"),
        (previous => "0100000110100100", load => '1', i => "0100001101000100", sel => "010101100", o => "0100001101000100"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "1101000011000101", sel => "001011111", o => "UUUUUUUUUUUUUUUU"),
        (previous => "0101011111110101", load => '0', i => "1101011110011010", sel => "001100001", o => "0101011111110101"),
        (previous => "0010010010011111", load => '0', i => "0000101100101001", sel => "011000001", o => "0010010010011111"),
        (previous => "0011001100001110", load => '0', i => "1011111101101110", sel => "011010100", o => "0011001100001110"),
        (previous => "1001000001101000", load => '1', i => "1111110000110111", sel => "000100000", o => "1111110000110111"),
        (previous => "1101000010110100", load => '0', i => "1010000010100100", sel => "011010011", o => "1101000010110100"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "1111011011111100", sel => "000010010", o => "1111011011111100"),
        (previous => "0010100110000111", load => '1', i => "0001101110110001", sel => "010111110", o => "0001101110110001"),
        (previous => "0001110111111101", load => '1', i => "0011001101011010", sel => "000100111", o => "0011001101011010"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "0100000000000110", sel => "010011011", o => "0100000000000110"),
        (previous => "1110000100110000", load => '0', i => "0001111001100101", sel => "011001010", o => "1110000100110000"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "1001001011000110", sel => "011010101", o => "1001001011000110"),
        (previous => "1100010001001111", load => '0', i => "0111011010001000", sel => "000100001", o => "1100010001001111"),
        (previous => "1000011110110110", load => '0', i => "1001111101011100", sel => "000110001", o => "1000011110110110"),
        (previous => "1010000011011000", load => '1', i => "1110110101111101", sel => "010011111", o => "1110110101111101"),
        (previous => "1101100101011101", load => '1', i => "0001101001010000", sel => "001100110", o => "0001101001010000"),
        (previous => "0111100001000000", load => '1', i => "1011110001100010", sel => "000101110", o => "1011110001100010"),
        (previous => "1101111100001100", load => '0', i => "0000001100100001", sel => "001001011", o => "1101111100001100"),
        (previous => "1100101011100000", load => '0', i => "0001001001001000", sel => "001011011", o => "1100101011100000"),
        (previous => "1001011010001101", load => '0', i => "1100100011100011", sel => "010101000", o => "1001011010001101"),
        (previous => "0000010100101111", load => '1', i => "1011101110101110", sel => "000111001", o => "1011101110101110"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "1000010110000011", sel => "010001111", o => "1000010110000011"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "1011101110100100", sel => "010000000", o => "1011101110100100"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "0110010011010101", sel => "010011010", o => "UUUUUUUUUUUUUUUU"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "0101111101110100", sel => "000100010", o => "0101111101110100"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "1011110011011011", sel => "011100001", o => "1011110011011011"),
        (previous => "1111001101100111", load => '1', i => "1100000100001001", sel => "001000100", o => "1100000100001001"),
        (previous => "0100010011000110", load => '0', i => "0000000001010101", sel => "010100011", o => "0100010011000110"),
        (previous => "0110001000000111", load => '0', i => "0001001110110000", sel => "010110011", o => "0110001000000111"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "1000100101011000", sel => "000011101", o => "UUUUUUUUUUUUUUUU"),
        (previous => "1000001011010111", load => '0', i => "1010010010010001", sel => "010001101", o => "1000001011010111"),
        (previous => "0011101110110011", load => '1', i => "0011011000100000", sel => "001100010", o => "0011011000100000"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "0001010110100001", sel => "011111110", o => "0001010110100001"),
        (previous => "1100010001001111", load => '0', i => "0100111000111011", sel => "000100001", o => "1100010001001111"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "1001111101011110", sel => "010100001", o => "UUUUUUUUUUUUUUUU"),
        (previous => "0100101011011000", load => '1', i => "0000010100111111", sel => "010011110", o => "0000010100111111"),
        (previous => "0011101000000000", load => '1', i => "0010000010000100", sel => "011101011", o => "0010000010000100"),
        (previous => "0100000000000110", load => '0', i => "1110100000100111", sel => "010011011", o => "0100000000000110"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "0111011111011011", sel => "001101011", o => "UUUUUUUUUUUUUUUU"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "0000001011111000", sel => "010000100", o => "UUUUUUUUUUUUUUUU"),
        (previous => "1011101110100100", load => '1', i => "1100100110000110", sel => "010000000", o => "1100100110000110"),
        (previous => "0101111010010100", load => '1', i => "1110100111101000", sel => "000101010", o => "1110100111101000"),
        (previous => "0011001001000111", load => '0', i => "1111011011100110", sel => "001010111", o => "0011001001000111"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "0110011100001000", sel => "000101000", o => "UUUUUUUUUUUUUUUU"),
        (previous => "0010011001111100", load => '0', i => "1101100110101001", sel => "011001110", o => "0010011001111100"),
        (previous => "0110010101110000", load => '1', i => "0011110001001000", sel => "011101000", o => "0011110001001000"),
        (previous => "0101101010001000", load => '1', i => "1010100100110011", sel => "011011110", o => "1010100100110011"),
        (previous => "0011010001001100", load => '1', i => "1101110011001110", sel => "011011101", o => "1101110011001110"),
        (previous => "1000011110110110", load => '0', i => "1101101000111010", sel => "000110001", o => "1000011110110110"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "1011001110111110", sel => "000110101", o => "UUUUUUUUUUUUUUUU"),
        (previous => "0111101100110010", load => '0', i => "0011001000111110", sel => "010010001", o => "0111101100110010"),
        (previous => "1110101111000011", load => '1', i => "0001000101101000", sel => "001111110", o => "0001000101101000"),
        (previous => "0110101101101010", load => '1', i => "1101011010111111", sel => "010001011", o => "1101011010111111"),
        (previous => "1110001111000001", load => '1', i => "0011110111100111", sel => "000111010", o => "0011110111100111"),
        (previous => "0010011011101001", load => '1', i => "1010101110110101", sel => "000100100", o => "1010101110110101"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "0111111110011101", sel => "001101100", o => "0111111110011101"),
        (previous => "0000000001000010", load => '0', i => "0111011001111011", sel => "011110011", o => "0000000001000010"),
        (previous => "1000011101100000", load => '1', i => "0101000101011000", sel => "011111111", o => "0101000101011000"),
        (previous => "0111010011001000", load => '1', i => "0001000010001001", sel => "000110010", o => "0001000010001001"),
        (previous => "1100001100101011", load => '1', i => "1100011110111110", sel => "001000000", o => "1100011110111110"),
        (previous => "1000001111011101", load => '1', i => "0000000001001111", sel => "001000110", o => "0000000001001111"),
        (previous => "1101000010110100", load => '1', i => "0101111011001101", sel => "011010011", o => "0101111011001101"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "0001100101011001", sel => "001001000", o => "UUUUUUUUUUUUUUUU"),
        (previous => "0100010011000110", load => '1', i => "0100010110010011", sel => "010100011", o => "0100010110010011"),
        (previous => "0000110100101111", load => '0', i => "0011000110110111", sel => "000000111", o => "0000110100101111"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "0111110100100011", sel => "000010100", o => "0111110100100011"),
        (previous => "0000001110010101", load => '1', i => "0010110100010110", sel => "001101001", o => "0010110100010110"),
        (previous => "0001000110001011", load => '1', i => "0110001000010101", sel => "011110001", o => "0110001000010101"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "0000010001000111", sel => "001001000", o => "0000010001000111"),
        (previous => "1000101111000111", load => '1', i => "1000101110000111", sel => "011011001", o => "1000101110000111"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "1111101011001110", sel => "000101000", o => "1111101011001110"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "0001101110100001", sel => "010110101", o => "UUUUUUUUUUUUUUUU"),
        (previous => "0011001101011111", load => '1', i => "1101011111101001", sel => "010101010", o => "1101011111101001"),
        (previous => "1011100100010011", load => '0', i => "0010011010001100", sel => "001011110", o => "1011100100010011"),
        (previous => "0011101011000000", load => '1', i => "0110111010010011", sel => "011111001", o => "0110111010010011"),
        (previous => "1101111000011111", load => '0', i => "1000100110100111", sel => "001001001", o => "1101111000011111"),
        (previous => "1001001010100011", load => '1', i => "1011010000010000", sel => "000110111", o => "1011010000010000"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "1001011100000010", sel => "010100000", o => "UUUUUUUUUUUUUUUU"),
        (previous => "0101011111110101", load => '0', i => "0000111101001010", sel => "001100001", o => "0101011111110101"),
        (previous => "0100001101000100", load => '1', i => "1111011100100100", sel => "010101100", o => "1111011100100100"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "0000001001001100", sel => "010110110", o => "0000001001001100"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "0110001100000010", sel => "000001111", o => "UUUUUUUUUUUUUUUU"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "0010101010101100", sel => "000110101", o => "0010101010101100"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "0011000000001011", sel => "010110101", o => "UUUUUUUUUUUUUUUU"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "1011000100000100", sel => "011000111", o => "1011000100000100"),
        (previous => "0111101100110010", load => '1', i => "0101100101001110", sel => "010010001", o => "0101100101001110"),
        (previous => "1100101000100011", load => '1', i => "1010100010000101", sel => "001111101", o => "1010100010000101"),
        (previous => "1100100110000110", load => '1', i => "0001010100100101", sel => "010000000", o => "0001010100100101"),
        (previous => "1011011111001011", load => '0', i => "1111000010000110", sel => "010011001", o => "1011011111001011"),
        (previous => "0110111010010011", load => '0', i => "0100101100110011", sel => "011111001", o => "0110111010010011"),
        (previous => "1010011000100110", load => '0', i => "1110110011101001", sel => "011100000", o => "1010011000100110"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "1101010111111000", sel => "010010110", o => "UUUUUUUUUUUUUUUU"),
        (previous => "0000001001111110", load => '1', i => "0110010100101101", sel => "011101100", o => "0110010100101101"),
        (previous => "0100100011011000", load => '0', i => "1011001111100010", sel => "000101100", o => "0100100011011000"),
        (previous => "0000010010010010", load => '0', i => "0000011110101010", sel => "011111000", o => "0000010010010010"),
        (previous => "0011001001000111", load => '0', i => "1001001000111011", sel => "001010111", o => "0011001001000111"),
        (previous => "1011100100010011", load => '1', i => "1101000010111000", sel => "001011110", o => "1101000010111000"),
        (previous => "0001101111101101", load => '0', i => "1111000000111001", sel => "001110110", o => "0001101111101101"),
        (previous => "1000010110000011", load => '1', i => "0101001011010010", sel => "010001111", o => "0101001011010010"),
        (previous => "0000000001000010", load => '0', i => "1111110011001011", sel => "011110011", o => "0000000001000010"),
        (previous => "0110010010000101", load => '1', i => "0111100110101011", sel => "001111011", o => "0111100110101011"),
        (previous => "0010010010010111", load => '1', i => "1100010001000001", sel => "001010000", o => "1100010001000001"),
        (previous => "0100101001000111", load => '0', i => "1111100000101110", sel => "000100110", o => "0100101001000111"),
        (previous => "0000010011011000", load => '1', i => "1110110101011010", sel => "010101001", o => "1110110101011010"),
        (previous => "1011010000010000", load => '1', i => "1100101001010010", sel => "000110111", o => "1100101001010010"),
        (previous => "1110000100110000", load => '0', i => "1111110110101001", sel => "011001010", o => "1110000100110000"),
        (previous => "1101011111101001", load => '0', i => "0001000100001000", sel => "010101010", o => "1101011111101001"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "1011100001111110", sel => "000010000", o => "1011100001111110"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "1000101100001101", sel => "010011010", o => "1000101100001101"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "1001100000000001", sel => "010101011", o => "UUUUUUUUUUUUUUUU"),
        (previous => "0101111001001011", load => '0', i => "1101011001111100", sel => "011101111", o => "0101111001001011"),
        (previous => "0010011011101111", load => '1', i => "0100100011001100", sel => "000011100", o => "0100100011001100"),
        (previous => "1100010000111010", load => '1', i => "0101000111110011", sel => "001000001", o => "0101000111110011"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "0001110010011100", sel => "010010100", o => "0001110010011100"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "1101100011010100", sel => "011001001", o => "1101100011010100"),
        (previous => "1001011010001101", load => '1', i => "0011011110011110", sel => "010101000", o => "0011011110011110"),
        (previous => "1110001101111101", load => '1', i => "1001001001001000", sel => "011000010", o => "1001001001001000"),
        (previous => "0001110010011100", load => '1', i => "1001000101011000", sel => "010010100", o => "1001000101011000"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "0100100111110011", sel => "010100000", o => "UUUUUUUUUUUUUUUU"),
        (previous => "1010100010000101", load => '1', i => "1010110010011110", sel => "001111101", o => "1010110010011110"),
        (previous => "0100101001000111", load => '0', i => "0000010010001110", sel => "000100110", o => "0100101001000111"),
        (previous => "0111001100001110", load => '0', i => "0011111010101010", sel => "001111010", o => "0111001100001110"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "0011000011101100", sel => "000001111", o => "0011000011101100"),
        (previous => "0101111011001101", load => '0', i => "0100000010000000", sel => "011010011", o => "0101111011001101"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "0010000101001001", sel => "011110000", o => "UUUUUUUUUUUUUUUU"),
        (previous => "0111011011000101", load => '0', i => "1101101011110001", sel => "001100000", o => "0111011011000101"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "1111111110110011", sel => "001111001", o => "UUUUUUUUUUUUUUUU"),
        (previous => "1000101100001101", load => '1', i => "0110000001000111", sel => "010011010", o => "0110000001000111"),
        (previous => "1011101110101110", load => '0', i => "1110110011100111", sel => "000111001", o => "1011101110101110"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "1111100001100101", sel => "011100101", o => "UUUUUUUUUUUUUUUU"),
        (previous => "1111010100010001", load => '0', i => "0111111110001011", sel => "010010011", o => "1111010100010001"),
        (previous => "1011100001111101", load => '1', i => "1111110000000101", sel => "010111101", o => "1111110000000101"),
        (previous => "0110001000000111", load => '1', i => "0011001000010100", sel => "010110011", o => "0011001000010100"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "0001100111100111", sel => "010011101", o => "0001100111100111"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "1010000011011000", sel => "000100011", o => "UUUUUUUUUUUUUUUU"),
        (previous => "1010110010011110", load => '1', i => "1001000100111000", sel => "001111101", o => "1001000100111000"),
        (previous => "0011000100100011", load => '0', i => "1110100010110001", sel => "001110101", o => "0011000100100011"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "1011100001001011", sel => "010110101", o => "1011100001001011"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "1011100010000100", sel => "001001110", o => "1011100010000100"),
        (previous => "1000100010000010", load => '0', i => "0111010001101001", sel => "011011010", o => "1000100010000010"),
        (previous => "1011100111011001", load => '1', i => "1000001111111100", sel => "000000101", o => "1000001111111100"),
        (previous => "1111110000000101", load => '0', i => "1011110110111001", sel => "010111101", o => "1111110000000101"),
        (previous => "1111110000110111", load => '0', i => "0110101001101101", sel => "000100000", o => "1111110000110111"),
        (previous => "0010100111010111", load => '0', i => "1101110000001010", sel => "001101111", o => "0010100111010111"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "0010111100101101", sel => "000111110", o => "UUUUUUUUUUUUUUUU"),
        (previous => "0000001101111111", load => '0', i => "0011110010101010", sel => "001010110", o => "0000001101111111"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "0011110000011111", sel => "001011111", o => "0011110000011111"),
        (previous => "0110101100110111", load => '0', i => "1011111111010100", sel => "000011011", o => "0110101100110111"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "0101100100100011", sel => "000011111", o => "UUUUUUUUUUUUUUUU"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "0101000111111101", sel => "000001010", o => "0101000111111101"),
        (previous => "1100100101011000", load => '0', i => "0101011100000010", sel => "001011010", o => "1100100101011000"),
        (previous => "0010101010101100", load => '1', i => "0110110011000000", sel => "000110101", o => "0110110011000000"),
        (previous => "0101111101110111", load => '0', i => "1101000111100000", sel => "000010101", o => "0101111101110111"),
        (previous => "0010000101110010", load => '0', i => "1011011101010000", sel => "000001001", o => "0010000101110010"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "0101110110001110", sel => "011100101", o => "0101110110001110"),
        (previous => "1011011111001011", load => '1', i => "1110010111100101", sel => "010011001", o => "1110010111100101"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "0010101101000100", sel => "010000101", o => "UUUUUUUUUUUUUUUU"),
        (previous => "0101111101110100", load => '1', i => "0010110101100000", sel => "000100010", o => "0010110101100000"),
        (previous => "0101000111111101", load => '0', i => "0100110001111111", sel => "000001010", o => "0101000111111101"),
        (previous => "0001101111101101", load => '1', i => "0111010110001001", sel => "001110110", o => "0111010110001001"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "1010000011100011", sel => "001001100", o => "UUUUUUUUUUUUUUUU"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "0100111000011000", sel => "000011110", o => "UUUUUUUUUUUUUUUU"),
        (previous => "1110110101011010", load => '0', i => "0111100100101101", sel => "010101001", o => "1110110101011010"),
        (previous => "1011110010111010", load => '0', i => "0101010000110110", sel => "010100010", o => "1011110010111010"),
        (previous => "0111111010001000", load => '1', i => "1111100100011100", sel => "010100100", o => "1111100100011100"),
        (previous => "0011001100001110", load => '0', i => "0000100010110101", sel => "011010100", o => "0011001100001110"),
        (previous => "0001110000000101", load => '0', i => "0001010000111011", sel => "010101101", o => "0001110000000101"),
        (previous => "0110111101011100", load => '0', i => "0000010001011101", sel => "010100110", o => "0110111101011100"),
        (previous => "0111111110101000", load => '1', i => "1001000101101000", sel => "001110011", o => "1001000101101000"),
        (previous => "1011111110111111", load => '0', i => "0111001111011110", sel => "001100011", o => "1011111110111111"),
        (previous => "1100010001000001", load => '1', i => "0010000000101010", sel => "001010000", o => "0010000000101010"),
        (previous => "1100011110111110", load => '1', i => "0001101001001000", sel => "001000000", o => "0001101001001000"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "0001111111110010", sel => "011110000", o => "UUUUUUUUUUUUUUUU"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "1001101110010100", sel => "010000001", o => "1001101110010100"),
        (previous => "0101011111110101", load => '1', i => "0110100100111000", sel => "001100001", o => "0110100100111000"),
        (previous => "1111010101000111", load => '0', i => "1011100000001100", sel => "011010000", o => "1111010101000111"),
        (previous => "1010101110110101", load => '1', i => "1100010010111010", sel => "000100100", o => "1100010010111010"),
        (previous => "1111110000000101", load => '1', i => "1100101101100000", sel => "010111101", o => "1100101101100000"),
        (previous => "1011100001001011", load => '1', i => "1000101111010011", sel => "010110101", o => "1000101111010011"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "0101111100110110", sel => "000101101", o => "0101111100110110"),
        (previous => "0101111100110110", load => '0', i => "1001011110000110", sel => "000101101", o => "0101111100110110"),
        (previous => "0101100110110010", load => '0', i => "1000101111000111", sel => "000010001", o => "0101100110110010"),
        (previous => "1000000110110111", load => '0', i => "1010100010110111", sel => "000001100", o => "1000000110110111"),
        (previous => "0110110011000000", load => '0', i => "1100000000111000", sel => "000110101", o => "0110110011000000"),
        (previous => "1001000101011000", load => '1', i => "1000100110011010", sel => "010010100", o => "1000100110011010"),
        (previous => "0011000011101100", load => '1', i => "0110001001101010", sel => "000001111", o => "0110001001101010"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "0011000010001111", sel => "000111111", o => "0011000010001111"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "0001111101001100", sel => "010101011", o => "0001111101001100"),
        (previous => "0010010101011100", load => '0', i => "0101110000000001", sel => "001110100", o => "0010010101011100"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "0011001100101110", sel => "010100101", o => "UUUUUUUUUUUUUUUU"),
        (previous => "0000111111010101", load => '1', i => "0001101001011100", sel => "010110100", o => "0001101001011100"),
        (previous => "0101001110000111", load => '0', i => "1011001001101101", sel => "011101110", o => "0101001110000111"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "0100100101111001", sel => "001110001", o => "0100100101111001"),
        (previous => "0101110110001110", load => '0', i => "0101100010101110", sel => "011100101", o => "0101110110001110"),
        (previous => "0101001110000111", load => '0', i => "0011010001000010", sel => "011101110", o => "0101001110000111"),
        (previous => "0000111001111000", load => '0', i => "1101010101010001", sel => "000101111", o => "0000111001111000"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "0100010010010001", sel => "001111100", o => "0100010010010001"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "1001011000111100", sel => "010000100", o => "1001011000111100"),
        (previous => "0010000010000100", load => '1', i => "1100111010110000", sel => "011101011", o => "1100111010110000"),
        (previous => "0100101001000111", load => '1', i => "0111111101010101", sel => "000100110", o => "0111111101010101"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "0001110000001001", sel => "010010110", o => "0001110000001001"),
        (previous => "1000001011010111", load => '0', i => "1100010011111000", sel => "010001101", o => "1000001011010111"),
        (previous => "1101111100001100", load => '0', i => "1001010001101001", sel => "001001011", o => "1101111100001100"),
        (previous => "0010010010011111", load => '0', i => "1010101001001110", sel => "011000001", o => "0010010010011111"),
        (previous => "0010100111010111", load => '1', i => "1010001000111100", sel => "001101111", o => "1010001000111100"),
        (previous => "1110101101010010", load => '0', i => "1110010101101011", sel => "010110111", o => "1110101101010010"),
        (previous => "0010110100010110", load => '1', i => "0010101111101000", sel => "001101001", o => "0010101111101000"),
        (previous => "0001111101001100", load => '1', i => "0011101001101100", sel => "010101011", o => "0011101001101100"),
        (previous => "0001100110101010", load => '1', i => "1101110001010111", sel => "000111000", o => "1101110001010111"),
        (previous => "1011000100000100", load => '0', i => "1001110101111101", sel => "011000111", o => "1011000100000100"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "1101110100010100", sel => "010000101", o => "UUUUUUUUUUUUUUUU"),
        (previous => "0000010100111111", load => '0', i => "0011001010100001", sel => "010011110", o => "0000010100111111"),
        (previous => "0011110001100100", load => '1', i => "0010100111101101", sel => "000100101", o => "0010100111101101"),
        (previous => "0010100111101101", load => '1', i => "0110101110101110", sel => "000100101", o => "0110101110101110"),
        (previous => "0101111011001101", load => '0', i => "1011100000011101", sel => "011010011", o => "0101111011001101"),
        (previous => "1110100001000111", load => '1', i => "1001100011010100", sel => "011000100", o => "1001100011010100"),
        (previous => "0000110100101111", load => '1', i => "0111000000111101", sel => "000000111", o => "0111000000111101"),
        (previous => "1000100010000010", load => '1', i => "0110111011101000", sel => "011011010", o => "0110111011101000"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "1011010000100001", sel => "011101010", o => "1011010000100001"),
        (previous => "1110110101011010", load => '0', i => "1001101111101000", sel => "010101001", o => "1110110101011010"),
        (previous => "0001101110110001", load => '0', i => "0101100101101101", sel => "010111110", o => "0001101110110001"),
        (previous => "0101011110000111", load => '0', i => "0000011100001100", sel => "011011100", o => "0101011110000111"),
        (previous => "0000111000110010", load => '1', i => "0101011100110001", sel => "011110010", o => "0101011100110001"),
        (previous => "0100100101111001", load => '1', i => "1001001101010110", sel => "001110001", o => "1001001101010110"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "0001010000101001", sel => "000111110", o => "UUUUUUUUUUUUUUUU"),
        (previous => "0000010001000111", load => '0', i => "0000110111101110", sel => "001001000", o => "0000010001000111"),
        (previous => "0001101110110001", load => '1', i => "0101010111110101", sel => "010111110", o => "0101010111110101"),
        (previous => "0110101100110111", load => '0', i => "0011000011001111", sel => "000011011", o => "0110101100110111"),
        (previous => "0101110110001110", load => '1', i => "0011010010111001", sel => "011100101", o => "0011010010111001"),
        (previous => "1001010010111010", load => '1', i => "0011000001100011", sel => "000000110", o => "0011000001100011"),
        (previous => "1111100100011100", load => '1', i => "1010001100100001", sel => "010100100", o => "1010001100100001"),
        (previous => "0011001001000111", load => '1', i => "1010100011111101", sel => "001010111", o => "1010100011111101"),
        (previous => "0011101001101100", load => '0', i => "0000011011101111", sel => "010101011", o => "0011101001101100"),
        (previous => "0110010100101101", load => '0', i => "0101000101100000", sel => "011101100", o => "0110010100101101"),
        (previous => "0010111011111110", load => '1', i => "0011001010011110", sel => "011011011", o => "0011001010011110"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "0100110011100111", sel => "011100111", o => "0100110011100111"),
        (previous => "1011000100000100", load => '0', i => "1000010110100101", sel => "011000111", o => "1011000100000100"),
        (previous => "0000110001011000", load => '0', i => "0000100011000000", sel => "011100100", o => "0000110001011000"),
        (previous => "1011010000100001", load => '1', i => "0001000010100101", sel => "011101010", o => "0001000010100101"),
        (previous => "0101100110110010", load => '0', i => "0111100110101011", sel => "000010001", o => "0101100110110010"),
        (previous => "1100010001001111", load => '1', i => "1110000101010000", sel => "000100001", o => "1110000101010000"),
        (previous => "0000010100111111", load => '0', i => "0010010010100111", sel => "010011110", o => "0000010100111111"),
        (previous => "0011001101011010", load => '1', i => "0111011001010010", sel => "000100111", o => "0111011001010010"),
        (previous => "1011110011011011", load => '1', i => "0000000000111110", sel => "011100001", o => "0000000000111110"),
        (previous => "0110001000010101", load => '0', i => "0010111000011001", sel => "011110001", o => "0110001000010101"),
        (previous => "1110100111101000", load => '1', i => "1011100000000000", sel => "000101010", o => "1011100000000000"),
        (previous => "1010010001001111", load => '0', i => "0011011011000111", sel => "001010010", o => "1010010001001111"),
        (previous => "1101001100101111", load => '0', i => "0001101010101011", sel => "001101110", o => "1101001100101111"),
        (previous => "1100100101011000", load => '0', i => "1101001010010110", sel => "001011010", o => "1100100101011000"),
        (previous => "0110001000110010", load => '1', i => "0001001010100111", sel => "000000000", o => "0001001010100111"),
        (previous => "0101110001111011", load => '1', i => "0111011011001000", sel => "000001000", o => "0111011011001000"),
        (previous => "0001000010001001", load => '0', i => "0101100001100110", sel => "000110010", o => "0001000010001001"),
        (previous => "1011100011010010", load => '0', i => "1011111010001101", sel => "001011000", o => "1011100011010010"),
        (previous => "1101001100101111", load => '0', i => "0000000001101110", sel => "001101110", o => "1101001100101111"),
        (previous => "1010101010000101", load => '1', i => "1011000101011111", sel => "011100011", o => "1011000101011111"),
        (previous => "1100111011110110", load => '1', i => "1110010110001010", sel => "011110111", o => "1110010110001010"),
        (previous => "0101011100110001", load => '0', i => "1010101011011100", sel => "011110010", o => "0101011100110001"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "0101011101001010", sel => "010010010", o => "UUUUUUUUUUUUUUUU"),
        (previous => "0000000001000010", load => '0', i => "0001101110100101", sel => "011110011", o => "0000000001000010"),
        (previous => "0110111010010011", load => '1', i => "0010110010100101", sel => "011111001", o => "0010110010100101"),
        (previous => "1101011111101001", load => '0', i => "1011101010101101", sel => "010101010", o => "1101011111101001"),
        (previous => "1111011100100100", load => '0', i => "0110100011011111", sel => "010101100", o => "1111011100100100"),
        (previous => "0010111101101100", load => '0', i => "1110000000111000", sel => "001010100", o => "0010111101101100"),
        (previous => "0000001000001111", load => '0', i => "0010011110100110", sel => "001001111", o => "0000001000001111"),
        (previous => "0000101011001110", load => '0', i => "1001000010001001", sel => "010000111", o => "0000101011001110"),
        (previous => "1000101110000111", load => '0', i => "0100110110000001", sel => "011011001", o => "1000101110000111"),
        (previous => "1011100000000000", load => '0', i => "1010101101110011", sel => "000101010", o => "1011100000000000"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "0011000000000110", sel => "001000011", o => "UUUUUUUUUUUUUUUU"),
        (previous => "0111000000111101", load => '1', i => "1110001111111001", sel => "000000111", o => "1110001111111001"),
        (previous => "0110100100111000", load => '0', i => "1101011111110010", sel => "001100001", o => "0110100100111000"),
        (previous => "0011011000100000", load => '0', i => "1000010110011100", sel => "001100010", o => "0011011000100000"),
        (previous => "0100100011011000", load => '1', i => "1100111001001000", sel => "000101100", o => "1100111001001000"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "1101011010011101", sel => "001011101", o => "1101011010011101"),
        (previous => "0110101100110111", load => '1', i => "0001010011101100", sel => "000011011", o => "0001010011101100"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "1000100101110011", sel => "001000111", o => "1000100101110011"),
        (previous => "0101111011001101", load => '0', i => "0110001001001100", sel => "011010011", o => "0101111011001101"),
        (previous => "1111010111101011", load => '1', i => "0101011101110111", sel => "011101001", o => "0101011101110111"),
        (previous => "0011001010011110", load => '1', i => "1001111110111010", sel => "011011011", o => "1001111110111010"),
        (previous => "1011000010010110", load => '0', i => "0101010111000001", sel => "000011000", o => "1011000010010110"),
        (previous => "0010110010100101", load => '0', i => "0100110000100010", sel => "011111001", o => "0010110010100101"),
        (previous => "0001010100100101", load => '1', i => "1001010110000100", sel => "010000000", o => "1001010110000100"),
        (previous => "0001101001011100", load => '1', i => "1010100010110001", sel => "010110100", o => "1010100010110001"),
        (previous => "1011000100000100", load => '0', i => "1101111000001110", sel => "011000111", o => "1011000100000100"),
        (previous => "0110000000110011", load => '0', i => "1111010000101001", sel => "000010011", o => "0110000000110011"),
        (previous => "0011011001110100", load => '0', i => "1110101101110000", sel => "000000100", o => "0011011001110100"),
        (previous => "0100110010101000", load => '0', i => "0111010101000100", sel => "001111111", o => "0100110010101000"),
        (previous => "0111100110101011", load => '1', i => "0111011100101101", sel => "001111011", o => "0111011100101101"),
        (previous => "1100111010110000", load => '1', i => "1001110000001001", sel => "011101011", o => "1001110000001001"),
        (previous => "0111011011000101", load => '0', i => "0011101100100001", sel => "001100000", o => "0111011011000101"),
        (previous => "0010011010100010", load => '0', i => "0111000000011010", sel => "011001111", o => "0010011010100010"),
        (previous => "0000111001111000", load => '1', i => "0110011110011010", sel => "000101111", o => "0110011110011010"),
        (previous => "1100111001001000", load => '0', i => "1101110001001110", sel => "000101100", o => "1100111001001000"),
        (previous => "0001111011101100", load => '0', i => "0011011100010110", sel => "001110010", o => "0001111011101100"),
        (previous => "0010111101101100", load => '1', i => "0101100000101001", sel => "001010100", o => "0101100000101001"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "0110011100101101", sel => "000100011", o => "0110011100101101"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "1111010010101101", sel => "001100101", o => "1111010010101101"),
        (previous => "0000000001000010", load => '1', i => "0100111000101000", sel => "011110011", o => "0100111000101000"),
        (previous => "0010110010100101", load => '0', i => "0001111100010011", sel => "011111001", o => "0010110010100101"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "1001011101110100", sel => "010111000", o => "1001011101110100"),
        (previous => "1011101110101110", load => '1', i => "1001101101000011", sel => "000111001", o => "1001101101000011"),
        (previous => "1001111110111010", load => '0', i => "0000001001110010", sel => "011011011", o => "1001111110111010"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "0101001010011111", sel => "000000010", o => "UUUUUUUUUUUUUUUU"),
        (previous => "0110111011101000", load => '0', i => "0101101000010001", sel => "011011010", o => "0110111011101000"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "1110111101100101", sel => "011000000", o => "1110111101100101"),
        (previous => "0010011010100010", load => '1', i => "0010011110001000", sel => "011001111", o => "0010011110001000"),
        (previous => "0000001000001111", load => '0', i => "1000101111101101", sel => "001001111", o => "0000001000001111"),
        (previous => "1111011011111100", load => '0', i => "0111111011100001", sel => "000010010", o => "1111011011111100"),
        (previous => "1011111001010010", load => '0', i => "0101011111011010", sel => "000000011", o => "1011111001010010"),
        (previous => "0101001100110001", load => '0', i => "1011011010010010", sel => "011111101", o => "0101001100110001"),
        (previous => "1011000010010110", load => '1', i => "1111000011001011", sel => "000011000", o => "1111000011001011"),
        (previous => "1011100010000100", load => '1', i => "0101001010100111", sel => "001001110", o => "0101001010100111"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "0111000110101001", sel => "000011110", o => "UUUUUUUUUUUUUUUU"),
        (previous => "1101000000100111", load => '1', i => "1111011010000100", sel => "000111100", o => "1111011010000100"),
        (previous => "1001001101010110", load => '1', i => "1011111101000100", sel => "001110001", o => "1011111101000100"),
        (previous => "0010011001111100", load => '1', i => "1100000000010100", sel => "011001110", o => "1100000000010100"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "1110010001100011", sel => "001011001", o => "1110010001100011"),
        (previous => "0101100101001110", load => '0', i => "1010000101110101", sel => "010010001", o => "0101100101001110"),
        (previous => "0101011100110001", load => '0', i => "0110111001111001", sel => "011110010", o => "0101011100110001"),
        (previous => "0001101001010000", load => '0', i => "1110011101110110", sel => "001100110", o => "0001101001010000"),
        (previous => "0101001010100111", load => '0', i => "0100011110001111", sel => "001001110", o => "0101001010100111"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "1111111011011101", sel => "001111001", o => "1111111011011101"),
        (previous => "0111001001010110", load => '0', i => "0111010011111011", sel => "000010110", o => "0111001001010110"),
        (previous => "1100111111001111", load => '0', i => "1000011000110111", sel => "001010011", o => "1100111111001111"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "0110100110101000", sel => "010100000", o => "0110100110101000"),
        (previous => "1100111111001111", load => '1', i => "0111011101110111", sel => "001010011", o => "0111011101110111"),
        (previous => "0101001011010010", load => '0', i => "0001011011010000", sel => "010001111", o => "0101001011010010"),
        (previous => "1001011101110100", load => '1', i => "0011110001100010", sel => "010111000", o => "0011110001100010"),
        (previous => "1001001001001000", load => '0', i => "0011011001010100", sel => "011000010", o => "1001001001001000"),
        (previous => "0110111101011100", load => '1', i => "0010001110111010", sel => "010100110", o => "0010001110111010"),
        (previous => "0100100011001100", load => '0', i => "1001110000001000", sel => "000011100", o => "0100100011001100"),
        (previous => "1101000010111000", load => '1', i => "0011101010000001", sel => "001011110", o => "0011101010000001"),
        (previous => "1000100101110011", load => '0', i => "0000000110010111", sel => "001000111", o => "1000100101110011"),
        (previous => "0110111011101000", load => '1', i => "0100001111101010", sel => "011011010", o => "0100001111101010"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "0101101110001011", sel => "011110000", o => "UUUUUUUUUUUUUUUU"),
        (previous => "1101111100001100", load => '1', i => "0011011111011110", sel => "001001011", o => "0011011111011110"),
        (previous => "0011111000001010", load => '1', i => "0000000001101101", sel => "010111010", o => "0000000001101101"),
        (previous => "1001100000100100", load => '1', i => "0100000100100101", sel => "010001100", o => "0100000100100101"),
        (previous => "0011001100001110", load => '1', i => "0111100011100111", sel => "011010100", o => "0111100011100111"),
        (previous => "1000100110011010", load => '1', i => "1111111110001101", sel => "010010100", o => "1111111110001101"),
        (previous => "0011010101001110", load => '1', i => "1000101110101010", sel => "011001011", o => "1000101110101010"),
        (previous => "0101100101001110", load => '0', i => "0000111000001000", sel => "010010001", o => "0101100101001110"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "1101100101010000", sel => "000110100", o => "UUUUUUUUUUUUUUUU"),
        (previous => "1000001000110010", load => '0', i => "0101111100101010", sel => "011010010", o => "1000001000110010"),
        (previous => "0011011110011110", load => '1', i => "1001011000011010", sel => "010101000", o => "1001011000011010"),
        (previous => "0111111101010101", load => '0', i => "0011110101100110", sel => "000100110", o => "0111111101010101"),
        (previous => "0001010011101100", load => '1', i => "0001010100100000", sel => "000011011", o => "0001010100100000"),
        (previous => "1010011000100110", load => '1', i => "0000000110101101", sel => "011100000", o => "0000000110101101"),
        (previous => "0111011011001000", load => '0', i => "1010010010000001", sel => "000001000", o => "0111011011001000"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "0110110000010101", sel => "010000011", o => "UUUUUUUUUUUUUUUU"),
        (previous => "1010001100101011", load => '0', i => "0011111111100001", sel => "010111001", o => "1010001100101011"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "0110011101110010", sel => "011110110", o => "UUUUUUUUUUUUUUUU"),
        (previous => "1000101111010011", load => '0', i => "1110000110100111", sel => "010110101", o => "1000101111010011"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "0010001101111001", sel => "000001011", o => "UUUUUUUUUUUUUUUU"),
        (previous => "0011011111011110", load => '1', i => "1011001100100001", sel => "001001011", o => "1011001100100001"),
        (previous => "1011100111001101", load => '1', i => "1111101001000111", sel => "000010111", o => "1111101001000111"),
        (previous => "0010010010011111", load => '1', i => "0111000001100010", sel => "011000001", o => "0111000001100010"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "0010110001000011", sel => "011011000", o => "UUUUUUUUUUUUUUUU"),
        (previous => "0101111101110111", load => '1', i => "0110101001001011", sel => "000010101", o => "0110101001001011"),
        (previous => "0011110111100111", load => '1', i => "0110000011001110", sel => "000111010", o => "0110000011001110"),
        (previous => "0110010100101101", load => '0', i => "0011001110000111", sel => "011101100", o => "0110010100101101"),
        (previous => "0000010001000111", load => '0', i => "0111111001111110", sel => "001001000", o => "0000010001000111"),
        (previous => "1111011100100100", load => '1', i => "0111110000110011", sel => "010101100", o => "0111110000110011"),
        (previous => "0110100100111000", load => '1', i => "0010111000111110", sel => "001100001", o => "0010111000111110"),
        (previous => "0011000010001111", load => '0', i => "1101100010001001", sel => "000111111", o => "0011000010001111"),
        (previous => "1101110001010111", load => '0', i => "1101011010100000", sel => "000111000", o => "1101110001010111"),
        (previous => "0001110101101001", load => '0', i => "0110000001100001", sel => "010010111", o => "0001110101101001"),
        (previous => "1111101001000111", load => '1', i => "0111011000111010", sel => "000010111", o => "0111011000111010"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "0101100101001111", sel => "001000011", o => "UUUUUUUUUUUUUUUU"),
        (previous => "0110001000010101", load => '1', i => "1000001010001001", sel => "011110001", o => "1000001010001001"),
        (previous => "1010100010110001", load => '0', i => "1111000101110101", sel => "010110100", o => "1010100010110001"),
        (previous => "1011100011010010", load => '0', i => "0011000110111101", sel => "001011000", o => "1011100011010010"),
        (previous => "1101001100101111", load => '1', i => "0101000101101010", sel => "001101110", o => "0101000101101010"),
        (previous => "1100111001001000", load => '1', i => "0010100111001011", sel => "000101100", o => "0010100111001011"),
        (previous => "1011111110111111", load => '1', i => "0001101000001010", sel => "001100011", o => "0001101000001010"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "1011100001000011", sel => "010111011", o => "1011100001000011"),
        (previous => "1100101011100000", load => '1', i => "0100000111011010", sel => "001011011", o => "0100000111011010"),
        (previous => "0011101010000001", load => '1', i => "1100101111110001", sel => "001011110", o => "1100101111110001"),
        (previous => "0100010110010011", load => '0', i => "0101100000110101", sel => "010100011", o => "0100010110010011"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "1000101100100110", sel => "000110100", o => "UUUUUUUUUUUUUUUU"),
        (previous => "1111010100010001", load => '1', i => "1101000011011010", sel => "010010011", o => "1101000011011010"),
        (previous => "1111111011011101", load => '1', i => "0110100100110010", sel => "001111001", o => "0110100100110010"),
        (previous => "1010100100110011", load => '1', i => "1011101110100000", sel => "011011110", o => "1011101110100000"),
        (previous => "0011000100100011", load => '0', i => "1010100111001100", sel => "001110101", o => "0011000100100011"),
        (previous => "1011001100100001", load => '0', i => "0101011100101111", sel => "001001011", o => "1011001100100001"),
        (previous => "1101011111101001", load => '1', i => "0111011011101011", sel => "010101010", o => "0111011011101011"),
        (previous => "1110110101011010", load => '0', i => "0000001101000110", sel => "010101001", o => "1110110101011010"),
        (previous => "0101000111111101", load => '1', i => "0110110010100100", sel => "000001010", o => "0110110010100100"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "1101111101001000", sel => "010100101", o => "UUUUUUUUUUUUUUUU"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "1100010101111100", sel => "010010000", o => "UUUUUUUUUUUUUUUU"),
        (previous => "0011011001110100", load => '0', i => "1000000000001111", sel => "000000100", o => "0011011001110100"),
        (previous => "1010000000001000", load => '0', i => "0100001010001000", sel => "011101101", o => "1010000000001000"),
        (previous => "1111111110001101", load => '1', i => "1000101101100110", sel => "010010100", o => "1000101101100110"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "1101011011011100", sel => "010100101", o => "1101011011011100"),
        (previous => "1001101110010100", load => '1', i => "0101001100100111", sel => "010000001", o => "0101001100100111"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "1101100011010001", sel => "001101000", o => "UUUUUUUUUUUUUUUU"),
        (previous => "0101100101001110", load => '0', i => "0011111001111010", sel => "010010001", o => "0101100101001110"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "1110010010000101", sel => "010010101", o => "1110010010000101"),
        (previous => "1101011010111111", load => '1', i => "0100000100101010", sel => "010001011", o => "0100000100101010"),
        (previous => "1000101111010011", load => '1', i => "1010110110111010", sel => "010110101", o => "1010110110111010"),
        (previous => "0011000001100011", load => '0', i => "1010110010111110", sel => "000000110", o => "0011000001100011"),
        (previous => "0101100011010111", load => '0', i => "0010111110101100", sel => "000110000", o => "0101100011010111"),
        (previous => "1000001011010111", load => '1', i => "0110100001000000", sel => "010001101", o => "0110100001000000"),
        (previous => "1010111011001110", load => '1', i => "1010011111100110", sel => "010001010", o => "1010011111100110"),
        (previous => "0111011101110111", load => '0', i => "0001100001100111", sel => "001010011", o => "0111011101110111"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "1101001111001111", sel => "001001100", o => "1101001111001111"),
        (previous => "0101100011010111", load => '1', i => "1001001001100001", sel => "000110000", o => "1001001001100001"),
        (previous => "0100000111011010", load => '0', i => "1001010111110110", sel => "001011011", o => "0100000111011010"),
        (previous => "1011100000000000", load => '1', i => "1010101010000001", sel => "000101010", o => "1010101010000001"),
        (previous => "0101000111110011", load => '1', i => "0010100000110111", sel => "001000001", o => "0010100000110111"),
        (previous => "0111100011100111", load => '0', i => "1001101000111101", sel => "011010100", o => "0111100011100111"),
        (previous => "0111010110001001", load => '0', i => "1101000101101101", sel => "001110110", o => "0111010110001001"),
        (previous => "0110100110101000", load => '0', i => "0011011011111010", sel => "010100000", o => "0110100110101000"),
        (previous => "1000011110110110", load => '0', i => "1000011010000100", sel => "000110001", o => "1000011110110110"),
        (previous => "0000010100111111", load => '0', i => "0110100111011000", sel => "010011110", o => "0000010100111111"),
        (previous => "0001000010001001", load => '1', i => "0011100000100100", sel => "000110010", o => "0011100000100100"),
        (previous => "0001110101101001", load => '0', i => "0110100001010101", sel => "010010111", o => "0001110101101001"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "1111110110110000", sel => "001110111", o => "1111110110110000"),
        (previous => "1001111110111010", load => '0', i => "0110010011011010", sel => "011011011", o => "1001111110111010"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "0111110100011011", sel => "001101010", o => "0111110100011011"),
        (previous => "1010100010110001", load => '0', i => "0000101111101111", sel => "010110100", o => "1010100010110001"),
        (previous => "0110001000101000", load => '0', i => "1001000101100101", sel => "010111100", o => "0110001000101000"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "0101000000000101", sel => "001110000", o => "UUUUUUUUUUUUUUUU"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "1101001100110111", sel => "001100100", o => "1101001100110111"),
        (previous => "0011000010001111", load => '1', i => "1111000111010101", sel => "000111111", o => "1111000111010101"),
        (previous => "0101001100100111", load => '1', i => "1111111100001000", sel => "010000001", o => "1111111100001000"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "1101001110011111", sel => "010010010", o => "UUUUUUUUUUUUUUUU"),
        (previous => "1000001111111100", load => '0', i => "1010111000010110", sel => "000000101", o => "1000001111111100"),
        (previous => "0101000101101010", load => '0', i => "0111001011110010", sel => "001101110", o => "0101000101101010"),
        (previous => "1011100011010010", load => '1', i => "0110001101011100", sel => "001011000", o => "0110001101011100"),
        (previous => "0111001100001110", load => '0', i => "0010110100010000", sel => "001111010", o => "0111001100001110"),
        (previous => "UUUUUUUUUUUUUUUU", load => '1', i => "0111110011001100", sel => "011011000", o => "0111110011001100"),
        (previous => "1010001100100001", load => '1', i => "1000001000111100", sel => "010100100", o => "1000001000111100"),
        (previous => "UUUUUUUUUUUUUUUU", load => '0', i => "1010010110100001", sel => "001101011", o => "UUUUUUUUUUUUUUUU"),
        (previous => "0000001001001100", load => '1', i => "1000111011100000", sel => "010110110", o => "1000111011100000"),
        (previous => "1000101110000111", load => '1', i => "0101011001100001", sel => "011011001", o => "0101011001100001")
    );
    CONSTANT total_cycles : INTEGER := test_cases'LENGTH;
    FUNCTION slv_to_string (slv : STD_LOGIC_VECTOR) RETURN STRING IS
        VARIABLE str : STRING (slv'length DOWNTO 1) := (OTHERS => NUL);
    BEGIN
        FOR n IN slv'length DOWNTO 1 LOOP
            str(n) := STD_LOGIC'image(slv((n - 1)))(2);
        END LOOP;
        RETURN str;
    END FUNCTION;

BEGIN
    bench : my_ram512 PORT MAP(clk, load, i, sel, o_actual);

    PROCESS
    BEGIN
        FOR cycle IN 1 TO total_cycles LOOP
            clk <= '0';
            WAIT FOR clk_period / 2;

            clk <= '1';
            WAIT FOR clk_period / 2;
        END LOOP;
        WAIT;
    END PROCESS;

    PROCESS
    BEGIN
        FOR n IN test_cases'RANGE LOOP
            previous <= test_cases(n).previous;
            i <= test_cases(n).i;
            load <= test_cases(n).load;
            sel <= test_cases(n).sel;

            WAIT FOR clk_period / 2;
            o_expected <= test_cases(n).o;
            WAIT FOR clk_period / 4;

            ASSERT (o_actual = o_expected)
            REPORT "test failed for " &
                "previous = " & slv_to_string(previous) &
                ". load = " & STD_LOGIC'image(load) &
                ". i = " & slv_to_string(i) &
                ". sel = " & slv_to_string(sel) &
                ". expected o = " & slv_to_string(o_expected) &
                ", got " & slv_to_string(o_actual) SEVERITY error;
            WAIT FOR clk_period / 4;
        END LOOP;
        WAIT;

    END PROCESS;

END behavioral;